
module AH_LruArbiter_64 (req
,gnt_busy
,gnt);

input [63:0] req;
input [63:0] gnt_busy;
output [63:0] gnt;


req [63:0] req0_used_status;
req [63:0] req1_used_status;
req [63:0] req2_used_status;
req [63:0] req3_used_status;
req [63:0] req4_used_status;
req [63:0] req5_used_status;
req [63:0] req6_used_status;
req [63:0] req7_used_status;
req [63:0] req8_used_status;
req [63:0] req9_used_status;
req [63:0] req10_used_status;
req [63:0] req11_used_status;
req [63:0] req12_used_status;
req [63:0] req13_used_status;
req [63:0] req14_used_status;
req [63:0] req15_used_status;
req [63:0] req16_used_status;
req [63:0] req17_used_status;
req [63:0] req18_used_status;
req [63:0] req19_used_status;
req [63:0] req20_used_status;
req [63:0] req21_used_status;
req [63:0] req22_used_status;
req [63:0] req23_used_status;
req [63:0] req24_used_status;
req [63:0] req25_used_status;
req [63:0] req26_used_status;
req [63:0] req27_used_status;
req [63:0] req28_used_status;
req [63:0] req29_used_status;
req [63:0] req30_used_status;
req [63:0] req31_used_status;
req [63:0] req32_used_status;
req [63:0] req33_used_status;
req [63:0] req34_used_status;
req [63:0] req35_used_status;
req [63:0] req36_used_status;
req [63:0] req37_used_status;
req [63:0] req38_used_status;
req [63:0] req39_used_status;
req [63:0] req40_used_status;
req [63:0] req41_used_status;
req [63:0] req42_used_status;
req [63:0] req43_used_status;
req [63:0] req44_used_status;
req [63:0] req45_used_status;
req [63:0] req46_used_status;
req [63:0] req47_used_status;
req [63:0] req48_used_status;
req [63:0] req49_used_status;
req [63:0] req50_used_status;
req [63:0] req51_used_status;
req [63:0] req52_used_status;
req [63:0] req53_used_status;
req [63:0] req54_used_status;
req [63:0] req55_used_status;
req [63:0] req56_used_status;
req [63:0] req57_used_status;
req [63:0] req58_used_status;
req [63:0] req59_used_status;
req [63:0] req60_used_status;
req [63:0] req61_used_status;
req [63:0] req62_used_status;
req [63:0] req63_used_status;

always @(posedge clk, negedge rstn) begin
        if(~rstn) begin

	req0_used_status <= 64'd64;
	req1_used_status <= 64'd63;
	req2_used_status <= 64'd62;
	req3_used_status <= 64'd61;
	req4_used_status <= 64'd60;
	req5_used_status <= 64'd59;
	req6_used_status <= 64'd58;
	req7_used_status <= 64'd57;
	req8_used_status <= 64'd56;
	req9_used_status <= 64'd55;
	req10_used_status <= 64'd54;
	req11_used_status <= 64'd53;
	req12_used_status <= 64'd52;
	req13_used_status <= 64'd51;
	req14_used_status <= 64'd50;
	req15_used_status <= 64'd49;
	req16_used_status <= 64'd48;
	req17_used_status <= 64'd47;
	req18_used_status <= 64'd46;
	req19_used_status <= 64'd45;
	req20_used_status <= 64'd44;
	req21_used_status <= 64'd43;
	req22_used_status <= 64'd42;
	req23_used_status <= 64'd41;
	req24_used_status <= 64'd40;
	req25_used_status <= 64'd39;
	req26_used_status <= 64'd38;
	req27_used_status <= 64'd37;
	req28_used_status <= 64'd36;
	req29_used_status <= 64'd35;
	req30_used_status <= 64'd34;
	req31_used_status <= 64'd33;
	req32_used_status <= 64'd32;
	req33_used_status <= 64'd31;
	req34_used_status <= 64'd30;
	req35_used_status <= 64'd29;
	req36_used_status <= 64'd28;
	req37_used_status <= 64'd27;
	req38_used_status <= 64'd26;
	req39_used_status <= 64'd25;
	req40_used_status <= 64'd24;
	req41_used_status <= 64'd23;
	req42_used_status <= 64'd22;
	req43_used_status <= 64'd21;
	req44_used_status <= 64'd20;
	req45_used_status <= 64'd19;
	req46_used_status <= 64'd18;
	req47_used_status <= 64'd17;
	req48_used_status <= 64'd16;
	req49_used_status <= 64'd15;
	req50_used_status <= 64'd14;
	req51_used_status <= 64'd13;
	req52_used_status <= 64'd12;
	req53_used_status <= 64'd11;
	req54_used_status <= 64'd10;
	req55_used_status <= 64'd9;
	req56_used_status <= 64'd8;
	req57_used_status <= 64'd7;
	req58_used_status <= 64'd6;
	req59_used_status <= 64'd5;
	req60_used_status <= 64'd4;
	req61_used_status <= 64'd3;
	req62_used_status <= 64'd2;
	req63_used_status <= 64'd1;

        end
        else begin

	gnt_pre[63:0] = 64'd0
	req_int[63:0]= req[64:0] & {64{gnt_busy}};
	if(req[0]) begin
		gnt_pre[0] = (req0_used_status==64) ? 1'b1 |

	((req1 & (req1_used_status > req0_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req0_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req0_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req0_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req0_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req0_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req0_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req0_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req0_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req0_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req0_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req0_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req0_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req0_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req0_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req0_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req0_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req0_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req0_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req0_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req0_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req0_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req0_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req0_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req0_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req0_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req0_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req0_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req0_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req0_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req0_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req0_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req0_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req0_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req0_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req0_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req0_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req0_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req0_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req0_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req0_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req0_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req0_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req0_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req0_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req0_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req0_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req0_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req0_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req0_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req0_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req0_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req0_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req0_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req0_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req0_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req0_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req0_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req0_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req0_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req0_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req0_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req0_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[1]) begin
		gnt_pre[1] = (req1_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req1_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req1_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req1_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req1_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req1_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req1_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req1_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req1_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req1_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req1_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req1_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req1_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req1_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req1_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req1_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req1_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req1_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req1_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req1_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req1_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req1_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req1_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req1_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req1_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req1_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req1_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req1_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req1_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req1_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req1_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req1_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req1_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req1_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req1_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req1_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req1_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req1_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req1_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req1_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req1_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req1_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req1_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req1_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req1_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req1_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req1_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req1_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req1_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req1_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req1_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req1_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req1_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req1_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req1_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req1_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req1_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req1_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req1_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req1_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req1_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req1_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req1_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req1_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[2]) begin
		gnt_pre[2] = (req2_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req2_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req2_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req2_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req2_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req2_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req2_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req2_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req2_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req2_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req2_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req2_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req2_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req2_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req2_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req2_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req2_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req2_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req2_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req2_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req2_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req2_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req2_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req2_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req2_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req2_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req2_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req2_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req2_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req2_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req2_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req2_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req2_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req2_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req2_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req2_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req2_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req2_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req2_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req2_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req2_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req2_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req2_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req2_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req2_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req2_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req2_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req2_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req2_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req2_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req2_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req2_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req2_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req2_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req2_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req2_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req2_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req2_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req2_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req2_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req2_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req2_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req2_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req2_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[3]) begin
		gnt_pre[3] = (req3_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req3_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req3_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req3_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req3_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req3_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req3_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req3_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req3_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req3_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req3_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req3_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req3_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req3_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req3_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req3_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req3_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req3_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req3_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req3_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req3_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req3_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req3_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req3_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req3_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req3_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req3_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req3_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req3_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req3_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req3_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req3_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req3_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req3_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req3_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req3_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req3_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req3_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req3_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req3_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req3_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req3_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req3_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req3_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req3_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req3_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req3_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req3_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req3_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req3_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req3_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req3_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req3_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req3_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req3_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req3_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req3_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req3_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req3_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req3_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req3_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req3_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req3_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req3_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[4]) begin
		gnt_pre[4] = (req4_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req4_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req4_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req4_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req4_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req4_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req4_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req4_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req4_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req4_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req4_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req4_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req4_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req4_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req4_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req4_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req4_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req4_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req4_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req4_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req4_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req4_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req4_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req4_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req4_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req4_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req4_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req4_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req4_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req4_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req4_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req4_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req4_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req4_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req4_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req4_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req4_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req4_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req4_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req4_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req4_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req4_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req4_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req4_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req4_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req4_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req4_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req4_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req4_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req4_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req4_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req4_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req4_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req4_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req4_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req4_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req4_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req4_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req4_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req4_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req4_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req4_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req4_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req4_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[5]) begin
		gnt_pre[5] = (req5_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req5_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req5_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req5_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req5_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req5_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req5_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req5_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req5_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req5_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req5_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req5_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req5_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req5_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req5_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req5_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req5_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req5_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req5_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req5_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req5_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req5_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req5_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req5_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req5_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req5_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req5_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req5_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req5_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req5_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req5_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req5_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req5_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req5_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req5_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req5_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req5_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req5_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req5_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req5_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req5_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req5_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req5_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req5_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req5_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req5_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req5_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req5_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req5_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req5_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req5_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req5_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req5_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req5_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req5_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req5_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req5_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req5_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req5_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req5_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req5_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req5_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req5_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req5_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[6]) begin
		gnt_pre[6] = (req6_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req6_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req6_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req6_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req6_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req6_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req6_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req6_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req6_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req6_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req6_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req6_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req6_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req6_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req6_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req6_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req6_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req6_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req6_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req6_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req6_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req6_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req6_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req6_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req6_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req6_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req6_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req6_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req6_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req6_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req6_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req6_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req6_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req6_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req6_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req6_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req6_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req6_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req6_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req6_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req6_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req6_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req6_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req6_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req6_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req6_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req6_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req6_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req6_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req6_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req6_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req6_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req6_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req6_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req6_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req6_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req6_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req6_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req6_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req6_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req6_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req6_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req6_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req6_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[7]) begin
		gnt_pre[7] = (req7_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req7_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req7_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req7_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req7_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req7_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req7_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req7_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req7_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req7_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req7_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req7_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req7_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req7_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req7_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req7_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req7_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req7_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req7_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req7_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req7_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req7_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req7_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req7_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req7_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req7_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req7_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req7_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req7_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req7_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req7_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req7_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req7_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req7_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req7_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req7_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req7_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req7_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req7_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req7_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req7_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req7_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req7_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req7_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req7_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req7_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req7_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req7_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req7_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req7_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req7_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req7_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req7_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req7_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req7_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req7_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req7_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req7_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req7_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req7_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req7_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req7_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req7_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req7_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[8]) begin
		gnt_pre[8] = (req8_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req8_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req8_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req8_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req8_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req8_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req8_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req8_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req8_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req8_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req8_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req8_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req8_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req8_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req8_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req8_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req8_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req8_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req8_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req8_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req8_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req8_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req8_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req8_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req8_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req8_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req8_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req8_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req8_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req8_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req8_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req8_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req8_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req8_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req8_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req8_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req8_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req8_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req8_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req8_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req8_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req8_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req8_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req8_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req8_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req8_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req8_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req8_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req8_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req8_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req8_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req8_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req8_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req8_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req8_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req8_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req8_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req8_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req8_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req8_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req8_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req8_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req8_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req8_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[9]) begin
		gnt_pre[9] = (req9_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req9_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req9_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req9_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req9_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req9_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req9_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req9_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req9_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req9_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req9_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req9_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req9_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req9_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req9_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req9_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req9_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req9_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req9_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req9_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req9_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req9_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req9_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req9_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req9_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req9_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req9_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req9_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req9_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req9_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req9_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req9_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req9_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req9_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req9_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req9_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req9_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req9_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req9_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req9_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req9_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req9_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req9_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req9_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req9_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req9_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req9_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req9_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req9_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req9_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req9_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req9_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req9_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req9_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req9_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req9_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req9_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req9_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req9_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req9_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req9_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req9_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req9_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req9_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[10]) begin
		gnt_pre[10] = (req10_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req10_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req10_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req10_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req10_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req10_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req10_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req10_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req10_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req10_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req10_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req10_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req10_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req10_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req10_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req10_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req10_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req10_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req10_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req10_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req10_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req10_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req10_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req10_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req10_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req10_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req10_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req10_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req10_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req10_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req10_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req10_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req10_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req10_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req10_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req10_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req10_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req10_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req10_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req10_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req10_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req10_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req10_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req10_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req10_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req10_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req10_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req10_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req10_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req10_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req10_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req10_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req10_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req10_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req10_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req10_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req10_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req10_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req10_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req10_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req10_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req10_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req10_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req10_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[11]) begin
		gnt_pre[11] = (req11_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req11_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req11_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req11_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req11_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req11_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req11_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req11_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req11_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req11_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req11_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req11_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req11_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req11_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req11_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req11_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req11_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req11_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req11_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req11_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req11_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req11_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req11_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req11_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req11_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req11_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req11_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req11_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req11_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req11_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req11_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req11_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req11_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req11_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req11_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req11_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req11_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req11_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req11_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req11_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req11_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req11_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req11_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req11_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req11_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req11_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req11_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req11_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req11_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req11_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req11_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req11_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req11_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req11_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req11_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req11_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req11_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req11_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req11_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req11_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req11_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req11_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req11_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req11_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[12]) begin
		gnt_pre[12] = (req12_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req12_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req12_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req12_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req12_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req12_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req12_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req12_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req12_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req12_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req12_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req12_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req12_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req12_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req12_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req12_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req12_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req12_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req12_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req12_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req12_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req12_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req12_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req12_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req12_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req12_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req12_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req12_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req12_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req12_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req12_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req12_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req12_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req12_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req12_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req12_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req12_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req12_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req12_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req12_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req12_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req12_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req12_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req12_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req12_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req12_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req12_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req12_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req12_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req12_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req12_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req12_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req12_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req12_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req12_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req12_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req12_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req12_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req12_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req12_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req12_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req12_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req12_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req12_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[13]) begin
		gnt_pre[13] = (req13_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req13_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req13_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req13_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req13_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req13_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req13_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req13_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req13_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req13_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req13_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req13_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req13_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req13_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req13_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req13_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req13_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req13_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req13_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req13_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req13_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req13_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req13_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req13_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req13_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req13_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req13_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req13_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req13_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req13_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req13_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req13_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req13_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req13_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req13_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req13_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req13_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req13_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req13_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req13_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req13_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req13_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req13_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req13_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req13_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req13_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req13_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req13_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req13_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req13_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req13_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req13_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req13_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req13_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req13_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req13_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req13_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req13_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req13_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req13_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req13_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req13_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req13_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req13_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[14]) begin
		gnt_pre[14] = (req14_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req14_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req14_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req14_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req14_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req14_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req14_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req14_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req14_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req14_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req14_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req14_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req14_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req14_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req14_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req14_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req14_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req14_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req14_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req14_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req14_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req14_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req14_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req14_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req14_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req14_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req14_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req14_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req14_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req14_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req14_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req14_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req14_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req14_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req14_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req14_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req14_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req14_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req14_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req14_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req14_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req14_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req14_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req14_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req14_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req14_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req14_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req14_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req14_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req14_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req14_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req14_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req14_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req14_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req14_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req14_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req14_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req14_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req14_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req14_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req14_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req14_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req14_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req14_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[15]) begin
		gnt_pre[15] = (req15_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req15_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req15_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req15_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req15_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req15_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req15_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req15_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req15_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req15_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req15_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req15_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req15_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req15_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req15_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req15_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req15_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req15_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req15_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req15_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req15_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req15_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req15_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req15_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req15_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req15_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req15_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req15_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req15_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req15_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req15_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req15_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req15_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req15_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req15_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req15_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req15_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req15_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req15_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req15_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req15_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req15_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req15_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req15_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req15_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req15_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req15_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req15_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req15_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req15_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req15_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req15_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req15_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req15_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req15_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req15_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req15_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req15_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req15_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req15_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req15_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req15_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req15_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req15_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[16]) begin
		gnt_pre[16] = (req16_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req16_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req16_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req16_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req16_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req16_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req16_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req16_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req16_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req16_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req16_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req16_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req16_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req16_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req16_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req16_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req16_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req16_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req16_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req16_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req16_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req16_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req16_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req16_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req16_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req16_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req16_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req16_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req16_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req16_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req16_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req16_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req16_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req16_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req16_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req16_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req16_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req16_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req16_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req16_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req16_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req16_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req16_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req16_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req16_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req16_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req16_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req16_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req16_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req16_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req16_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req16_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req16_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req16_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req16_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req16_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req16_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req16_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req16_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req16_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req16_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req16_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req16_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req16_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[17]) begin
		gnt_pre[17] = (req17_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req17_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req17_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req17_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req17_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req17_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req17_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req17_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req17_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req17_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req17_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req17_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req17_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req17_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req17_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req17_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req17_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req17_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req17_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req17_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req17_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req17_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req17_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req17_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req17_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req17_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req17_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req17_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req17_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req17_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req17_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req17_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req17_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req17_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req17_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req17_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req17_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req17_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req17_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req17_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req17_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req17_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req17_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req17_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req17_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req17_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req17_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req17_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req17_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req17_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req17_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req17_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req17_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req17_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req17_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req17_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req17_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req17_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req17_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req17_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req17_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req17_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req17_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req17_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[18]) begin
		gnt_pre[18] = (req18_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req18_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req18_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req18_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req18_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req18_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req18_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req18_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req18_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req18_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req18_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req18_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req18_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req18_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req18_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req18_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req18_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req18_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req18_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req18_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req18_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req18_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req18_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req18_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req18_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req18_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req18_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req18_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req18_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req18_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req18_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req18_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req18_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req18_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req18_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req18_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req18_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req18_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req18_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req18_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req18_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req18_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req18_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req18_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req18_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req18_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req18_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req18_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req18_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req18_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req18_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req18_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req18_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req18_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req18_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req18_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req18_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req18_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req18_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req18_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req18_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req18_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req18_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req18_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[19]) begin
		gnt_pre[19] = (req19_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req19_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req19_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req19_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req19_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req19_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req19_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req19_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req19_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req19_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req19_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req19_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req19_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req19_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req19_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req19_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req19_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req19_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req19_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req19_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req19_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req19_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req19_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req19_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req19_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req19_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req19_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req19_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req19_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req19_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req19_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req19_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req19_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req19_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req19_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req19_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req19_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req19_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req19_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req19_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req19_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req19_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req19_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req19_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req19_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req19_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req19_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req19_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req19_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req19_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req19_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req19_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req19_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req19_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req19_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req19_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req19_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req19_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req19_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req19_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req19_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req19_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req19_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req19_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[20]) begin
		gnt_pre[20] = (req20_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req20_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req20_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req20_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req20_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req20_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req20_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req20_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req20_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req20_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req20_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req20_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req20_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req20_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req20_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req20_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req20_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req20_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req20_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req20_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req20_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req20_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req20_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req20_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req20_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req20_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req20_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req20_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req20_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req20_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req20_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req20_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req20_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req20_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req20_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req20_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req20_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req20_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req20_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req20_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req20_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req20_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req20_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req20_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req20_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req20_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req20_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req20_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req20_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req20_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req20_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req20_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req20_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req20_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req20_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req20_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req20_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req20_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req20_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req20_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req20_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req20_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req20_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req20_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[21]) begin
		gnt_pre[21] = (req21_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req21_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req21_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req21_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req21_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req21_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req21_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req21_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req21_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req21_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req21_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req21_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req21_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req21_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req21_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req21_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req21_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req21_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req21_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req21_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req21_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req21_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req21_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req21_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req21_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req21_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req21_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req21_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req21_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req21_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req21_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req21_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req21_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req21_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req21_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req21_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req21_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req21_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req21_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req21_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req21_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req21_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req21_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req21_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req21_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req21_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req21_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req21_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req21_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req21_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req21_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req21_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req21_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req21_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req21_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req21_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req21_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req21_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req21_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req21_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req21_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req21_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req21_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req21_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[22]) begin
		gnt_pre[22] = (req22_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req22_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req22_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req22_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req22_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req22_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req22_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req22_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req22_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req22_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req22_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req22_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req22_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req22_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req22_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req22_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req22_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req22_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req22_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req22_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req22_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req22_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req22_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req22_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req22_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req22_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req22_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req22_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req22_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req22_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req22_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req22_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req22_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req22_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req22_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req22_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req22_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req22_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req22_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req22_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req22_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req22_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req22_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req22_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req22_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req22_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req22_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req22_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req22_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req22_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req22_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req22_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req22_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req22_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req22_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req22_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req22_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req22_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req22_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req22_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req22_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req22_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req22_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req22_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[23]) begin
		gnt_pre[23] = (req23_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req23_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req23_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req23_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req23_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req23_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req23_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req23_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req23_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req23_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req23_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req23_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req23_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req23_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req23_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req23_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req23_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req23_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req23_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req23_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req23_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req23_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req23_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req23_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req23_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req23_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req23_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req23_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req23_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req23_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req23_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req23_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req23_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req23_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req23_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req23_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req23_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req23_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req23_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req23_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req23_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req23_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req23_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req23_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req23_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req23_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req23_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req23_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req23_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req23_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req23_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req23_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req23_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req23_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req23_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req23_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req23_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req23_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req23_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req23_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req23_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req23_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req23_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req23_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[24]) begin
		gnt_pre[24] = (req24_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req24_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req24_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req24_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req24_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req24_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req24_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req24_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req24_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req24_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req24_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req24_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req24_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req24_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req24_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req24_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req24_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req24_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req24_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req24_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req24_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req24_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req24_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req24_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req24_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req24_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req24_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req24_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req24_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req24_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req24_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req24_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req24_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req24_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req24_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req24_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req24_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req24_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req24_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req24_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req24_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req24_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req24_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req24_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req24_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req24_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req24_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req24_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req24_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req24_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req24_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req24_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req24_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req24_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req24_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req24_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req24_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req24_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req24_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req24_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req24_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req24_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req24_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req24_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[25]) begin
		gnt_pre[25] = (req25_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req25_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req25_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req25_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req25_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req25_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req25_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req25_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req25_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req25_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req25_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req25_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req25_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req25_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req25_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req25_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req25_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req25_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req25_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req25_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req25_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req25_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req25_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req25_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req25_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req25_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req25_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req25_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req25_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req25_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req25_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req25_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req25_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req25_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req25_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req25_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req25_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req25_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req25_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req25_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req25_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req25_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req25_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req25_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req25_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req25_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req25_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req25_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req25_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req25_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req25_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req25_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req25_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req25_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req25_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req25_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req25_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req25_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req25_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req25_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req25_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req25_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req25_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req25_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[26]) begin
		gnt_pre[26] = (req26_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req26_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req26_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req26_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req26_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req26_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req26_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req26_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req26_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req26_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req26_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req26_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req26_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req26_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req26_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req26_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req26_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req26_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req26_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req26_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req26_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req26_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req26_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req26_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req26_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req26_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req26_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req26_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req26_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req26_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req26_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req26_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req26_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req26_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req26_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req26_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req26_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req26_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req26_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req26_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req26_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req26_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req26_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req26_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req26_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req26_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req26_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req26_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req26_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req26_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req26_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req26_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req26_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req26_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req26_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req26_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req26_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req26_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req26_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req26_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req26_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req26_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req26_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req26_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[27]) begin
		gnt_pre[27] = (req27_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req27_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req27_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req27_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req27_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req27_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req27_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req27_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req27_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req27_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req27_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req27_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req27_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req27_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req27_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req27_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req27_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req27_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req27_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req27_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req27_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req27_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req27_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req27_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req27_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req27_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req27_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req27_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req27_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req27_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req27_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req27_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req27_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req27_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req27_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req27_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req27_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req27_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req27_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req27_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req27_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req27_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req27_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req27_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req27_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req27_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req27_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req27_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req27_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req27_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req27_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req27_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req27_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req27_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req27_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req27_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req27_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req27_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req27_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req27_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req27_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req27_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req27_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req27_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[28]) begin
		gnt_pre[28] = (req28_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req28_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req28_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req28_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req28_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req28_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req28_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req28_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req28_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req28_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req28_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req28_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req28_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req28_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req28_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req28_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req28_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req28_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req28_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req28_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req28_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req28_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req28_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req28_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req28_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req28_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req28_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req28_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req28_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req28_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req28_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req28_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req28_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req28_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req28_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req28_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req28_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req28_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req28_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req28_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req28_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req28_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req28_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req28_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req28_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req28_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req28_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req28_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req28_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req28_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req28_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req28_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req28_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req28_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req28_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req28_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req28_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req28_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req28_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req28_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req28_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req28_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req28_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req28_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[29]) begin
		gnt_pre[29] = (req29_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req29_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req29_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req29_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req29_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req29_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req29_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req29_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req29_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req29_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req29_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req29_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req29_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req29_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req29_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req29_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req29_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req29_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req29_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req29_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req29_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req29_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req29_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req29_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req29_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req29_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req29_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req29_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req29_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req29_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req29_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req29_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req29_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req29_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req29_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req29_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req29_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req29_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req29_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req29_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req29_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req29_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req29_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req29_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req29_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req29_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req29_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req29_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req29_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req29_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req29_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req29_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req29_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req29_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req29_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req29_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req29_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req29_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req29_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req29_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req29_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req29_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req29_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req29_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[30]) begin
		gnt_pre[30] = (req30_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req30_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req30_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req30_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req30_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req30_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req30_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req30_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req30_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req30_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req30_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req30_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req30_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req30_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req30_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req30_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req30_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req30_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req30_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req30_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req30_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req30_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req30_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req30_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req30_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req30_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req30_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req30_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req30_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req30_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req30_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req30_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req30_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req30_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req30_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req30_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req30_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req30_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req30_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req30_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req30_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req30_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req30_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req30_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req30_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req30_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req30_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req30_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req30_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req30_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req30_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req30_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req30_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req30_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req30_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req30_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req30_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req30_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req30_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req30_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req30_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req30_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req30_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req30_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[31]) begin
		gnt_pre[31] = (req31_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req31_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req31_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req31_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req31_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req31_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req31_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req31_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req31_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req31_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req31_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req31_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req31_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req31_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req31_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req31_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req31_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req31_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req31_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req31_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req31_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req31_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req31_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req31_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req31_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req31_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req31_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req31_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req31_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req31_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req31_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req31_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req31_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req31_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req31_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req31_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req31_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req31_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req31_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req31_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req31_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req31_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req31_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req31_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req31_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req31_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req31_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req31_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req31_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req31_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req31_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req31_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req31_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req31_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req31_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req31_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req31_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req31_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req31_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req31_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req31_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req31_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req31_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req31_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[32]) begin
		gnt_pre[32] = (req32_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req32_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req32_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req32_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req32_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req32_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req32_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req32_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req32_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req32_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req32_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req32_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req32_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req32_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req32_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req32_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req32_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req32_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req32_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req32_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req32_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req32_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req32_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req32_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req32_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req32_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req32_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req32_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req32_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req32_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req32_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req32_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req32_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req32_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req32_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req32_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req32_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req32_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req32_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req32_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req32_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req32_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req32_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req32_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req32_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req32_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req32_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req32_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req32_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req32_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req32_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req32_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req32_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req32_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req32_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req32_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req32_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req32_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req32_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req32_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req32_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req32_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req32_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req32_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[33]) begin
		gnt_pre[33] = (req33_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req33_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req33_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req33_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req33_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req33_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req33_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req33_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req33_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req33_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req33_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req33_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req33_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req33_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req33_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req33_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req33_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req33_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req33_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req33_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req33_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req33_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req33_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req33_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req33_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req33_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req33_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req33_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req33_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req33_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req33_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req33_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req33_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req33_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req33_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req33_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req33_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req33_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req33_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req33_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req33_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req33_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req33_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req33_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req33_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req33_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req33_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req33_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req33_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req33_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req33_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req33_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req33_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req33_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req33_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req33_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req33_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req33_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req33_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req33_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req33_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req33_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req33_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req33_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[34]) begin
		gnt_pre[34] = (req34_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req34_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req34_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req34_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req34_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req34_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req34_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req34_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req34_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req34_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req34_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req34_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req34_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req34_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req34_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req34_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req34_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req34_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req34_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req34_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req34_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req34_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req34_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req34_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req34_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req34_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req34_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req34_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req34_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req34_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req34_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req34_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req34_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req34_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req34_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req34_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req34_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req34_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req34_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req34_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req34_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req34_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req34_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req34_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req34_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req34_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req34_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req34_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req34_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req34_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req34_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req34_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req34_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req34_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req34_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req34_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req34_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req34_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req34_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req34_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req34_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req34_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req34_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req34_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[35]) begin
		gnt_pre[35] = (req35_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req35_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req35_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req35_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req35_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req35_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req35_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req35_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req35_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req35_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req35_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req35_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req35_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req35_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req35_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req35_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req35_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req35_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req35_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req35_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req35_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req35_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req35_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req35_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req35_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req35_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req35_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req35_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req35_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req35_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req35_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req35_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req35_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req35_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req35_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req35_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req35_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req35_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req35_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req35_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req35_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req35_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req35_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req35_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req35_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req35_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req35_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req35_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req35_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req35_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req35_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req35_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req35_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req35_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req35_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req35_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req35_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req35_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req35_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req35_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req35_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req35_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req35_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req35_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[36]) begin
		gnt_pre[36] = (req36_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req36_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req36_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req36_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req36_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req36_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req36_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req36_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req36_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req36_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req36_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req36_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req36_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req36_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req36_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req36_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req36_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req36_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req36_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req36_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req36_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req36_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req36_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req36_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req36_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req36_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req36_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req36_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req36_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req36_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req36_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req36_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req36_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req36_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req36_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req36_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req36_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req36_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req36_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req36_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req36_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req36_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req36_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req36_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req36_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req36_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req36_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req36_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req36_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req36_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req36_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req36_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req36_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req36_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req36_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req36_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req36_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req36_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req36_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req36_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req36_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req36_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req36_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req36_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[37]) begin
		gnt_pre[37] = (req37_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req37_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req37_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req37_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req37_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req37_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req37_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req37_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req37_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req37_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req37_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req37_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req37_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req37_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req37_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req37_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req37_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req37_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req37_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req37_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req37_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req37_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req37_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req37_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req37_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req37_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req37_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req37_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req37_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req37_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req37_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req37_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req37_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req37_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req37_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req37_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req37_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req37_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req37_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req37_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req37_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req37_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req37_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req37_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req37_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req37_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req37_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req37_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req37_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req37_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req37_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req37_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req37_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req37_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req37_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req37_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req37_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req37_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req37_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req37_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req37_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req37_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req37_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req37_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[38]) begin
		gnt_pre[38] = (req38_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req38_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req38_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req38_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req38_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req38_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req38_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req38_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req38_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req38_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req38_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req38_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req38_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req38_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req38_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req38_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req38_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req38_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req38_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req38_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req38_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req38_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req38_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req38_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req38_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req38_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req38_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req38_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req38_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req38_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req38_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req38_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req38_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req38_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req38_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req38_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req38_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req38_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req38_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req38_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req38_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req38_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req38_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req38_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req38_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req38_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req38_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req38_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req38_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req38_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req38_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req38_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req38_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req38_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req38_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req38_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req38_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req38_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req38_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req38_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req38_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req38_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req38_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req38_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[39]) begin
		gnt_pre[39] = (req39_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req39_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req39_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req39_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req39_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req39_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req39_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req39_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req39_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req39_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req39_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req39_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req39_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req39_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req39_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req39_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req39_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req39_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req39_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req39_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req39_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req39_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req39_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req39_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req39_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req39_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req39_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req39_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req39_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req39_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req39_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req39_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req39_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req39_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req39_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req39_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req39_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req39_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req39_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req39_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req39_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req39_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req39_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req39_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req39_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req39_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req39_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req39_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req39_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req39_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req39_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req39_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req39_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req39_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req39_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req39_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req39_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req39_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req39_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req39_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req39_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req39_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req39_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req39_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[40]) begin
		gnt_pre[40] = (req40_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req40_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req40_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req40_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req40_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req40_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req40_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req40_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req40_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req40_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req40_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req40_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req40_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req40_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req40_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req40_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req40_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req40_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req40_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req40_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req40_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req40_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req40_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req40_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req40_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req40_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req40_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req40_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req40_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req40_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req40_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req40_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req40_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req40_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req40_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req40_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req40_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req40_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req40_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req40_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req40_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req40_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req40_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req40_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req40_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req40_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req40_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req40_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req40_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req40_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req40_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req40_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req40_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req40_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req40_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req40_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req40_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req40_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req40_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req40_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req40_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req40_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req40_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req40_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[41]) begin
		gnt_pre[41] = (req41_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req41_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req41_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req41_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req41_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req41_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req41_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req41_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req41_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req41_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req41_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req41_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req41_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req41_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req41_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req41_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req41_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req41_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req41_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req41_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req41_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req41_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req41_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req41_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req41_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req41_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req41_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req41_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req41_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req41_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req41_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req41_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req41_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req41_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req41_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req41_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req41_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req41_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req41_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req41_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req41_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req41_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req41_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req41_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req41_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req41_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req41_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req41_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req41_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req41_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req41_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req41_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req41_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req41_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req41_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req41_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req41_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req41_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req41_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req41_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req41_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req41_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req41_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req41_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[42]) begin
		gnt_pre[42] = (req42_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req42_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req42_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req42_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req42_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req42_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req42_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req42_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req42_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req42_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req42_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req42_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req42_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req42_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req42_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req42_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req42_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req42_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req42_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req42_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req42_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req42_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req42_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req42_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req42_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req42_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req42_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req42_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req42_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req42_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req42_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req42_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req42_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req42_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req42_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req42_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req42_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req42_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req42_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req42_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req42_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req42_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req42_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req42_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req42_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req42_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req42_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req42_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req42_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req42_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req42_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req42_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req42_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req42_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req42_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req42_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req42_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req42_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req42_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req42_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req42_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req42_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req42_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req42_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[43]) begin
		gnt_pre[43] = (req43_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req43_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req43_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req43_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req43_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req43_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req43_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req43_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req43_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req43_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req43_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req43_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req43_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req43_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req43_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req43_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req43_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req43_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req43_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req43_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req43_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req43_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req43_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req43_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req43_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req43_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req43_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req43_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req43_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req43_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req43_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req43_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req43_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req43_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req43_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req43_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req43_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req43_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req43_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req43_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req43_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req43_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req43_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req43_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req43_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req43_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req43_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req43_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req43_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req43_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req43_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req43_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req43_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req43_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req43_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req43_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req43_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req43_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req43_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req43_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req43_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req43_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req43_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req43_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[44]) begin
		gnt_pre[44] = (req44_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req44_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req44_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req44_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req44_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req44_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req44_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req44_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req44_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req44_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req44_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req44_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req44_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req44_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req44_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req44_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req44_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req44_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req44_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req44_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req44_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req44_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req44_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req44_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req44_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req44_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req44_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req44_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req44_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req44_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req44_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req44_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req44_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req44_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req44_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req44_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req44_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req44_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req44_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req44_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req44_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req44_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req44_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req44_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req44_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req44_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req44_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req44_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req44_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req44_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req44_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req44_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req44_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req44_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req44_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req44_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req44_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req44_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req44_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req44_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req44_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req44_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req44_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req44_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[45]) begin
		gnt_pre[45] = (req45_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req45_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req45_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req45_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req45_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req45_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req45_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req45_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req45_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req45_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req45_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req45_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req45_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req45_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req45_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req45_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req45_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req45_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req45_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req45_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req45_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req45_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req45_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req45_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req45_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req45_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req45_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req45_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req45_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req45_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req45_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req45_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req45_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req45_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req45_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req45_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req45_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req45_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req45_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req45_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req45_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req45_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req45_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req45_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req45_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req45_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req45_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req45_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req45_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req45_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req45_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req45_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req45_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req45_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req45_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req45_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req45_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req45_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req45_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req45_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req45_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req45_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req45_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req45_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[46]) begin
		gnt_pre[46] = (req46_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req46_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req46_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req46_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req46_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req46_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req46_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req46_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req46_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req46_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req46_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req46_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req46_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req46_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req46_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req46_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req46_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req46_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req46_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req46_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req46_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req46_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req46_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req46_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req46_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req46_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req46_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req46_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req46_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req46_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req46_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req46_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req46_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req46_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req46_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req46_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req46_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req46_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req46_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req46_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req46_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req46_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req46_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req46_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req46_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req46_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req46_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req46_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req46_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req46_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req46_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req46_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req46_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req46_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req46_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req46_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req46_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req46_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req46_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req46_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req46_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req46_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req46_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req46_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[47]) begin
		gnt_pre[47] = (req47_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req47_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req47_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req47_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req47_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req47_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req47_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req47_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req47_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req47_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req47_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req47_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req47_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req47_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req47_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req47_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req47_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req47_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req47_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req47_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req47_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req47_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req47_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req47_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req47_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req47_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req47_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req47_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req47_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req47_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req47_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req47_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req47_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req47_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req47_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req47_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req47_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req47_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req47_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req47_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req47_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req47_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req47_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req47_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req47_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req47_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req47_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req47_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req47_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req47_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req47_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req47_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req47_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req47_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req47_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req47_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req47_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req47_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req47_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req47_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req47_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req47_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req47_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req47_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[48]) begin
		gnt_pre[48] = (req48_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req48_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req48_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req48_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req48_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req48_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req48_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req48_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req48_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req48_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req48_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req48_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req48_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req48_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req48_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req48_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req48_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req48_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req48_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req48_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req48_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req48_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req48_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req48_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req48_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req48_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req48_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req48_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req48_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req48_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req48_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req48_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req48_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req48_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req48_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req48_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req48_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req48_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req48_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req48_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req48_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req48_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req48_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req48_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req48_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req48_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req48_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req48_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req48_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req48_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req48_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req48_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req48_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req48_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req48_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req48_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req48_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req48_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req48_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req48_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req48_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req48_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req48_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req48_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[49]) begin
		gnt_pre[49] = (req49_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req49_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req49_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req49_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req49_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req49_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req49_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req49_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req49_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req49_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req49_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req49_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req49_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req49_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req49_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req49_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req49_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req49_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req49_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req49_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req49_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req49_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req49_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req49_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req49_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req49_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req49_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req49_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req49_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req49_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req49_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req49_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req49_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req49_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req49_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req49_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req49_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req49_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req49_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req49_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req49_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req49_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req49_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req49_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req49_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req49_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req49_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req49_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req49_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req49_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req49_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req49_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req49_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req49_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req49_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req49_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req49_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req49_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req49_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req49_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req49_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req49_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req49_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req49_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[50]) begin
		gnt_pre[50] = (req50_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req50_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req50_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req50_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req50_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req50_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req50_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req50_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req50_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req50_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req50_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req50_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req50_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req50_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req50_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req50_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req50_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req50_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req50_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req50_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req50_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req50_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req50_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req50_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req50_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req50_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req50_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req50_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req50_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req50_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req50_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req50_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req50_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req50_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req50_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req50_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req50_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req50_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req50_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req50_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req50_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req50_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req50_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req50_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req50_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req50_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req50_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req50_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req50_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req50_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req50_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req50_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req50_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req50_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req50_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req50_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req50_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req50_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req50_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req50_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req50_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req50_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req50_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req50_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[51]) begin
		gnt_pre[51] = (req51_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req51_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req51_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req51_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req51_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req51_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req51_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req51_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req51_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req51_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req51_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req51_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req51_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req51_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req51_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req51_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req51_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req51_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req51_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req51_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req51_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req51_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req51_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req51_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req51_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req51_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req51_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req51_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req51_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req51_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req51_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req51_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req51_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req51_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req51_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req51_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req51_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req51_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req51_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req51_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req51_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req51_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req51_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req51_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req51_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req51_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req51_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req51_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req51_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req51_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req51_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req51_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req51_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req51_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req51_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req51_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req51_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req51_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req51_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req51_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req51_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req51_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req51_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req51_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[52]) begin
		gnt_pre[52] = (req52_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req52_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req52_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req52_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req52_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req52_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req52_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req52_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req52_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req52_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req52_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req52_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req52_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req52_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req52_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req52_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req52_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req52_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req52_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req52_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req52_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req52_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req52_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req52_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req52_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req52_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req52_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req52_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req52_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req52_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req52_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req52_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req52_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req52_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req52_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req52_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req52_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req52_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req52_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req52_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req52_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req52_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req52_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req52_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req52_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req52_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req52_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req52_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req52_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req52_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req52_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req52_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req52_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req52_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req52_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req52_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req52_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req52_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req52_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req52_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req52_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req52_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req52_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req52_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[53]) begin
		gnt_pre[53] = (req53_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req53_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req53_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req53_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req53_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req53_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req53_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req53_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req53_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req53_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req53_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req53_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req53_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req53_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req53_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req53_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req53_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req53_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req53_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req53_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req53_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req53_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req53_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req53_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req53_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req53_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req53_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req53_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req53_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req53_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req53_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req53_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req53_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req53_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req53_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req53_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req53_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req53_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req53_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req53_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req53_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req53_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req53_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req53_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req53_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req53_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req53_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req53_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req53_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req53_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req53_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req53_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req53_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req53_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req53_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req53_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req53_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req53_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req53_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req53_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req53_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req53_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req53_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req53_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[54]) begin
		gnt_pre[54] = (req54_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req54_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req54_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req54_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req54_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req54_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req54_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req54_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req54_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req54_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req54_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req54_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req54_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req54_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req54_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req54_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req54_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req54_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req54_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req54_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req54_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req54_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req54_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req54_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req54_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req54_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req54_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req54_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req54_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req54_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req54_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req54_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req54_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req54_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req54_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req54_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req54_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req54_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req54_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req54_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req54_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req54_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req54_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req54_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req54_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req54_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req54_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req54_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req54_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req54_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req54_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req54_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req54_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req54_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req54_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req54_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req54_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req54_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req54_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req54_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req54_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req54_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req54_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req54_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[55]) begin
		gnt_pre[55] = (req55_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req55_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req55_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req55_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req55_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req55_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req55_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req55_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req55_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req55_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req55_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req55_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req55_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req55_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req55_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req55_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req55_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req55_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req55_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req55_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req55_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req55_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req55_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req55_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req55_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req55_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req55_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req55_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req55_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req55_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req55_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req55_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req55_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req55_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req55_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req55_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req55_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req55_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req55_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req55_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req55_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req55_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req55_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req55_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req55_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req55_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req55_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req55_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req55_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req55_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req55_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req55_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req55_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req55_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req55_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req55_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req55_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req55_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req55_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req55_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req55_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req55_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req55_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req55_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[56]) begin
		gnt_pre[56] = (req56_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req56_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req56_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req56_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req56_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req56_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req56_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req56_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req56_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req56_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req56_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req56_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req56_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req56_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req56_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req56_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req56_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req56_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req56_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req56_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req56_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req56_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req56_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req56_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req56_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req56_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req56_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req56_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req56_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req56_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req56_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req56_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req56_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req56_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req56_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req56_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req56_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req56_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req56_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req56_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req56_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req56_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req56_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req56_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req56_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req56_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req56_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req56_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req56_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req56_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req56_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req56_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req56_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req56_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req56_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req56_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req56_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req56_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req56_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req56_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req56_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req56_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req56_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req56_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[57]) begin
		gnt_pre[57] = (req57_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req57_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req57_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req57_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req57_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req57_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req57_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req57_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req57_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req57_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req57_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req57_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req57_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req57_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req57_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req57_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req57_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req57_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req57_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req57_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req57_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req57_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req57_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req57_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req57_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req57_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req57_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req57_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req57_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req57_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req57_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req57_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req57_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req57_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req57_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req57_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req57_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req57_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req57_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req57_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req57_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req57_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req57_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req57_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req57_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req57_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req57_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req57_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req57_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req57_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req57_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req57_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req57_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req57_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req57_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req57_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req57_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req57_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req57_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req57_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req57_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req57_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req57_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req57_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[58]) begin
		gnt_pre[58] = (req58_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req58_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req58_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req58_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req58_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req58_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req58_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req58_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req58_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req58_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req58_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req58_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req58_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req58_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req58_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req58_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req58_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req58_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req58_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req58_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req58_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req58_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req58_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req58_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req58_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req58_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req58_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req58_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req58_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req58_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req58_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req58_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req58_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req58_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req58_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req58_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req58_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req58_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req58_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req58_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req58_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req58_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req58_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req58_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req58_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req58_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req58_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req58_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req58_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req58_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req58_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req58_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req58_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req58_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req58_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req58_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req58_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req58_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req58_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req58_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req58_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req58_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req58_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req58_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[59]) begin
		gnt_pre[59] = (req59_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req59_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req59_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req59_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req59_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req59_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req59_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req59_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req59_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req59_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req59_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req59_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req59_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req59_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req59_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req59_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req59_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req59_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req59_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req59_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req59_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req59_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req59_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req59_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req59_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req59_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req59_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req59_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req59_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req59_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req59_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req59_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req59_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req59_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req59_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req59_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req59_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req59_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req59_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req59_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req59_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req59_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req59_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req59_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req59_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req59_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req59_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req59_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req59_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req59_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req59_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req59_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req59_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req59_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req59_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req59_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req59_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req59_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req59_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req59_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req59_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req59_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req59_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req59_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[60]) begin
		gnt_pre[60] = (req60_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req60_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req60_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req60_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req60_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req60_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req60_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req60_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req60_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req60_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req60_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req60_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req60_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req60_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req60_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req60_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req60_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req60_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req60_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req60_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req60_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req60_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req60_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req60_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req60_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req60_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req60_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req60_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req60_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req60_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req60_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req60_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req60_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req60_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req60_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req60_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req60_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req60_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req60_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req60_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req60_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req60_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req60_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req60_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req60_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req60_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req60_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req60_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req60_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req60_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req60_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req60_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req60_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req60_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req60_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req60_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req60_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req60_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req60_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req60_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req60_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req60_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req60_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req60_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[61]) begin
		gnt_pre[61] = (req61_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req61_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req61_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req61_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req61_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req61_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req61_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req61_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req61_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req61_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req61_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req61_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req61_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req61_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req61_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req61_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req61_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req61_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req61_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req61_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req61_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req61_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req61_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req61_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req61_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req61_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req61_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req61_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req61_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req61_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req61_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req61_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req61_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req61_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req61_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req61_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req61_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req61_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req61_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req61_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req61_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req61_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req61_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req61_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req61_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req61_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req61_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req61_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req61_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req61_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req61_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req61_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req61_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req61_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req61_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req61_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req61_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req61_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req61_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req61_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req61_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req61_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req61_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req61_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[62]) begin
		gnt_pre[62] = (req62_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req62_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req62_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req62_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req62_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req62_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req62_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req62_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req62_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req62_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req62_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req62_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req62_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req62_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req62_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req62_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req62_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req62_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req62_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req62_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req62_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req62_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req62_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req62_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req62_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req62_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req62_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req62_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req62_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req62_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req62_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req62_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req62_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req62_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req62_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req62_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req62_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req62_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req62_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req62_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req62_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req62_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req62_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req62_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req62_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req62_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req62_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req62_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req62_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req62_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req62_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req62_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req62_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req62_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req62_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req62_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req62_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req62_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req62_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req62_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req62_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req62_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req62_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req62_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[63]) begin
		gnt_pre[63] = (req63_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req63_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req63_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req63_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req63_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req63_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req63_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req63_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req63_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req63_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req63_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req63_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req63_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req63_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req63_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req63_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req63_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req63_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req63_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req63_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req63_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req63_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req63_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req63_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req63_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req63_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req63_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req63_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req63_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req63_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req63_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req63_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req63_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req63_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req63_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req63_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req63_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req63_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req63_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req63_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req63_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req63_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req63_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req63_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req63_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req63_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req63_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req63_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req63_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req63_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req63_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req63_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req63_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req63_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req63_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req63_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req63_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req63_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req63_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req63_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req63_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req63_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req63_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req63_used_status)) ?1'b0 |
		1'b1;
	end

always @(req, gnt_busy) begin

	gnt_pre[63:0] = 64'd0
	req_int[63:0]= req[64:0] & {64{gnt_busy}};
	if(req[0]) begin
		gnt_pre[0] = (req0_used_status==64) ? 1'b1 |

	((req1 & (req1_used_status > req0_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req0_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req0_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req0_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req0_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req0_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req0_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req0_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req0_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req0_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req0_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req0_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req0_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req0_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req0_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req0_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req0_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req0_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req0_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req0_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req0_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req0_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req0_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req0_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req0_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req0_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req0_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req0_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req0_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req0_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req0_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req0_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req0_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req0_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req0_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req0_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req0_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req0_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req0_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req0_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req0_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req0_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req0_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req0_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req0_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req0_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req0_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req0_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req0_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req0_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req0_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req0_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req0_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req0_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req0_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req0_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req0_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req0_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req0_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req0_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req0_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req0_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req0_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[1]) begin
		gnt_pre[1] = (req1_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req1_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req1_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req1_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req1_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req1_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req1_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req1_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req1_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req1_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req1_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req1_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req1_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req1_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req1_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req1_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req1_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req1_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req1_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req1_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req1_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req1_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req1_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req1_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req1_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req1_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req1_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req1_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req1_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req1_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req1_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req1_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req1_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req1_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req1_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req1_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req1_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req1_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req1_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req1_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req1_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req1_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req1_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req1_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req1_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req1_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req1_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req1_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req1_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req1_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req1_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req1_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req1_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req1_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req1_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req1_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req1_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req1_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req1_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req1_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req1_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req1_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req1_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req1_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[2]) begin
		gnt_pre[2] = (req2_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req2_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req2_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req2_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req2_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req2_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req2_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req2_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req2_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req2_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req2_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req2_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req2_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req2_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req2_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req2_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req2_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req2_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req2_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req2_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req2_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req2_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req2_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req2_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req2_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req2_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req2_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req2_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req2_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req2_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req2_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req2_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req2_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req2_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req2_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req2_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req2_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req2_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req2_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req2_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req2_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req2_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req2_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req2_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req2_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req2_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req2_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req2_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req2_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req2_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req2_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req2_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req2_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req2_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req2_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req2_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req2_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req2_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req2_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req2_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req2_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req2_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req2_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req2_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[3]) begin
		gnt_pre[3] = (req3_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req3_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req3_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req3_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req3_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req3_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req3_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req3_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req3_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req3_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req3_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req3_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req3_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req3_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req3_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req3_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req3_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req3_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req3_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req3_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req3_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req3_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req3_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req3_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req3_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req3_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req3_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req3_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req3_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req3_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req3_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req3_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req3_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req3_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req3_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req3_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req3_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req3_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req3_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req3_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req3_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req3_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req3_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req3_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req3_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req3_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req3_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req3_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req3_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req3_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req3_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req3_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req3_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req3_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req3_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req3_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req3_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req3_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req3_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req3_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req3_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req3_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req3_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req3_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[4]) begin
		gnt_pre[4] = (req4_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req4_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req4_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req4_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req4_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req4_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req4_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req4_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req4_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req4_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req4_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req4_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req4_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req4_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req4_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req4_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req4_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req4_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req4_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req4_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req4_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req4_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req4_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req4_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req4_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req4_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req4_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req4_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req4_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req4_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req4_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req4_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req4_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req4_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req4_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req4_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req4_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req4_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req4_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req4_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req4_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req4_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req4_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req4_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req4_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req4_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req4_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req4_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req4_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req4_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req4_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req4_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req4_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req4_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req4_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req4_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req4_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req4_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req4_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req4_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req4_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req4_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req4_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req4_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[5]) begin
		gnt_pre[5] = (req5_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req5_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req5_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req5_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req5_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req5_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req5_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req5_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req5_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req5_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req5_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req5_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req5_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req5_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req5_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req5_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req5_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req5_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req5_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req5_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req5_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req5_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req5_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req5_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req5_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req5_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req5_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req5_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req5_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req5_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req5_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req5_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req5_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req5_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req5_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req5_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req5_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req5_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req5_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req5_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req5_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req5_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req5_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req5_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req5_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req5_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req5_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req5_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req5_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req5_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req5_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req5_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req5_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req5_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req5_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req5_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req5_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req5_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req5_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req5_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req5_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req5_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req5_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req5_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[6]) begin
		gnt_pre[6] = (req6_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req6_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req6_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req6_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req6_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req6_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req6_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req6_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req6_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req6_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req6_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req6_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req6_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req6_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req6_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req6_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req6_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req6_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req6_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req6_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req6_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req6_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req6_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req6_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req6_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req6_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req6_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req6_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req6_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req6_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req6_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req6_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req6_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req6_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req6_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req6_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req6_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req6_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req6_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req6_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req6_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req6_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req6_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req6_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req6_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req6_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req6_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req6_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req6_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req6_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req6_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req6_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req6_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req6_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req6_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req6_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req6_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req6_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req6_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req6_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req6_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req6_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req6_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req6_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[7]) begin
		gnt_pre[7] = (req7_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req7_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req7_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req7_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req7_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req7_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req7_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req7_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req7_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req7_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req7_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req7_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req7_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req7_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req7_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req7_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req7_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req7_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req7_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req7_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req7_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req7_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req7_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req7_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req7_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req7_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req7_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req7_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req7_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req7_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req7_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req7_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req7_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req7_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req7_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req7_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req7_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req7_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req7_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req7_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req7_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req7_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req7_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req7_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req7_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req7_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req7_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req7_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req7_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req7_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req7_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req7_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req7_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req7_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req7_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req7_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req7_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req7_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req7_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req7_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req7_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req7_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req7_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req7_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[8]) begin
		gnt_pre[8] = (req8_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req8_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req8_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req8_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req8_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req8_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req8_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req8_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req8_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req8_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req8_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req8_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req8_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req8_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req8_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req8_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req8_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req8_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req8_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req8_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req8_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req8_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req8_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req8_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req8_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req8_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req8_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req8_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req8_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req8_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req8_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req8_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req8_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req8_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req8_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req8_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req8_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req8_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req8_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req8_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req8_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req8_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req8_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req8_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req8_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req8_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req8_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req8_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req8_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req8_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req8_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req8_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req8_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req8_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req8_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req8_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req8_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req8_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req8_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req8_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req8_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req8_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req8_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req8_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[9]) begin
		gnt_pre[9] = (req9_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req9_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req9_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req9_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req9_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req9_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req9_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req9_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req9_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req9_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req9_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req9_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req9_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req9_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req9_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req9_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req9_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req9_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req9_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req9_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req9_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req9_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req9_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req9_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req9_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req9_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req9_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req9_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req9_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req9_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req9_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req9_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req9_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req9_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req9_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req9_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req9_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req9_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req9_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req9_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req9_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req9_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req9_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req9_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req9_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req9_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req9_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req9_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req9_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req9_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req9_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req9_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req9_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req9_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req9_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req9_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req9_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req9_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req9_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req9_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req9_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req9_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req9_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req9_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[10]) begin
		gnt_pre[10] = (req10_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req10_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req10_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req10_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req10_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req10_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req10_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req10_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req10_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req10_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req10_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req10_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req10_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req10_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req10_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req10_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req10_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req10_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req10_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req10_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req10_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req10_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req10_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req10_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req10_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req10_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req10_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req10_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req10_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req10_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req10_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req10_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req10_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req10_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req10_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req10_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req10_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req10_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req10_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req10_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req10_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req10_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req10_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req10_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req10_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req10_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req10_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req10_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req10_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req10_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req10_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req10_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req10_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req10_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req10_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req10_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req10_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req10_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req10_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req10_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req10_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req10_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req10_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req10_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[11]) begin
		gnt_pre[11] = (req11_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req11_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req11_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req11_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req11_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req11_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req11_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req11_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req11_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req11_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req11_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req11_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req11_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req11_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req11_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req11_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req11_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req11_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req11_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req11_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req11_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req11_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req11_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req11_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req11_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req11_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req11_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req11_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req11_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req11_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req11_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req11_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req11_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req11_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req11_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req11_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req11_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req11_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req11_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req11_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req11_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req11_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req11_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req11_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req11_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req11_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req11_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req11_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req11_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req11_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req11_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req11_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req11_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req11_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req11_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req11_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req11_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req11_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req11_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req11_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req11_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req11_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req11_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req11_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[12]) begin
		gnt_pre[12] = (req12_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req12_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req12_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req12_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req12_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req12_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req12_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req12_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req12_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req12_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req12_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req12_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req12_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req12_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req12_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req12_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req12_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req12_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req12_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req12_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req12_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req12_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req12_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req12_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req12_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req12_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req12_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req12_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req12_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req12_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req12_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req12_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req12_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req12_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req12_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req12_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req12_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req12_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req12_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req12_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req12_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req12_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req12_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req12_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req12_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req12_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req12_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req12_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req12_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req12_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req12_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req12_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req12_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req12_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req12_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req12_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req12_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req12_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req12_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req12_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req12_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req12_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req12_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req12_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[13]) begin
		gnt_pre[13] = (req13_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req13_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req13_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req13_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req13_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req13_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req13_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req13_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req13_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req13_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req13_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req13_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req13_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req13_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req13_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req13_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req13_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req13_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req13_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req13_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req13_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req13_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req13_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req13_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req13_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req13_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req13_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req13_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req13_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req13_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req13_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req13_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req13_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req13_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req13_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req13_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req13_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req13_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req13_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req13_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req13_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req13_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req13_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req13_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req13_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req13_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req13_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req13_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req13_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req13_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req13_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req13_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req13_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req13_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req13_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req13_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req13_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req13_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req13_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req13_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req13_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req13_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req13_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req13_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[14]) begin
		gnt_pre[14] = (req14_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req14_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req14_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req14_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req14_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req14_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req14_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req14_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req14_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req14_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req14_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req14_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req14_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req14_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req14_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req14_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req14_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req14_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req14_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req14_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req14_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req14_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req14_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req14_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req14_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req14_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req14_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req14_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req14_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req14_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req14_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req14_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req14_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req14_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req14_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req14_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req14_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req14_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req14_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req14_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req14_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req14_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req14_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req14_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req14_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req14_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req14_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req14_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req14_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req14_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req14_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req14_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req14_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req14_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req14_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req14_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req14_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req14_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req14_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req14_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req14_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req14_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req14_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req14_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[15]) begin
		gnt_pre[15] = (req15_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req15_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req15_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req15_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req15_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req15_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req15_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req15_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req15_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req15_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req15_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req15_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req15_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req15_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req15_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req15_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req15_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req15_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req15_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req15_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req15_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req15_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req15_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req15_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req15_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req15_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req15_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req15_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req15_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req15_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req15_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req15_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req15_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req15_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req15_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req15_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req15_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req15_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req15_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req15_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req15_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req15_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req15_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req15_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req15_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req15_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req15_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req15_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req15_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req15_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req15_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req15_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req15_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req15_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req15_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req15_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req15_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req15_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req15_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req15_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req15_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req15_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req15_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req15_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[16]) begin
		gnt_pre[16] = (req16_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req16_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req16_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req16_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req16_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req16_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req16_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req16_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req16_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req16_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req16_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req16_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req16_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req16_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req16_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req16_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req16_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req16_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req16_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req16_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req16_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req16_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req16_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req16_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req16_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req16_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req16_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req16_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req16_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req16_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req16_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req16_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req16_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req16_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req16_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req16_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req16_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req16_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req16_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req16_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req16_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req16_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req16_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req16_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req16_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req16_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req16_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req16_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req16_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req16_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req16_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req16_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req16_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req16_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req16_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req16_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req16_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req16_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req16_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req16_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req16_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req16_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req16_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req16_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[17]) begin
		gnt_pre[17] = (req17_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req17_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req17_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req17_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req17_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req17_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req17_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req17_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req17_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req17_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req17_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req17_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req17_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req17_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req17_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req17_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req17_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req17_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req17_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req17_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req17_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req17_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req17_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req17_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req17_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req17_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req17_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req17_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req17_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req17_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req17_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req17_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req17_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req17_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req17_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req17_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req17_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req17_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req17_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req17_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req17_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req17_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req17_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req17_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req17_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req17_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req17_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req17_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req17_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req17_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req17_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req17_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req17_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req17_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req17_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req17_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req17_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req17_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req17_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req17_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req17_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req17_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req17_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req17_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[18]) begin
		gnt_pre[18] = (req18_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req18_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req18_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req18_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req18_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req18_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req18_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req18_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req18_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req18_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req18_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req18_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req18_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req18_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req18_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req18_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req18_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req18_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req18_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req18_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req18_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req18_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req18_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req18_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req18_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req18_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req18_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req18_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req18_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req18_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req18_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req18_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req18_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req18_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req18_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req18_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req18_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req18_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req18_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req18_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req18_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req18_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req18_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req18_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req18_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req18_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req18_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req18_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req18_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req18_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req18_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req18_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req18_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req18_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req18_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req18_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req18_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req18_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req18_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req18_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req18_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req18_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req18_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req18_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[19]) begin
		gnt_pre[19] = (req19_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req19_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req19_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req19_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req19_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req19_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req19_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req19_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req19_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req19_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req19_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req19_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req19_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req19_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req19_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req19_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req19_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req19_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req19_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req19_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req19_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req19_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req19_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req19_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req19_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req19_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req19_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req19_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req19_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req19_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req19_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req19_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req19_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req19_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req19_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req19_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req19_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req19_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req19_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req19_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req19_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req19_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req19_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req19_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req19_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req19_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req19_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req19_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req19_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req19_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req19_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req19_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req19_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req19_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req19_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req19_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req19_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req19_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req19_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req19_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req19_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req19_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req19_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req19_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[20]) begin
		gnt_pre[20] = (req20_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req20_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req20_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req20_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req20_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req20_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req20_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req20_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req20_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req20_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req20_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req20_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req20_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req20_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req20_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req20_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req20_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req20_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req20_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req20_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req20_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req20_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req20_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req20_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req20_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req20_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req20_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req20_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req20_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req20_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req20_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req20_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req20_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req20_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req20_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req20_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req20_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req20_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req20_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req20_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req20_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req20_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req20_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req20_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req20_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req20_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req20_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req20_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req20_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req20_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req20_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req20_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req20_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req20_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req20_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req20_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req20_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req20_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req20_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req20_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req20_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req20_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req20_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req20_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[21]) begin
		gnt_pre[21] = (req21_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req21_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req21_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req21_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req21_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req21_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req21_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req21_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req21_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req21_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req21_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req21_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req21_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req21_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req21_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req21_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req21_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req21_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req21_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req21_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req21_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req21_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req21_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req21_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req21_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req21_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req21_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req21_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req21_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req21_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req21_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req21_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req21_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req21_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req21_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req21_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req21_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req21_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req21_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req21_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req21_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req21_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req21_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req21_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req21_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req21_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req21_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req21_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req21_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req21_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req21_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req21_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req21_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req21_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req21_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req21_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req21_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req21_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req21_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req21_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req21_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req21_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req21_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req21_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[22]) begin
		gnt_pre[22] = (req22_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req22_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req22_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req22_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req22_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req22_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req22_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req22_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req22_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req22_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req22_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req22_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req22_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req22_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req22_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req22_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req22_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req22_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req22_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req22_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req22_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req22_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req22_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req22_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req22_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req22_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req22_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req22_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req22_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req22_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req22_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req22_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req22_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req22_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req22_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req22_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req22_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req22_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req22_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req22_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req22_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req22_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req22_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req22_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req22_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req22_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req22_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req22_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req22_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req22_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req22_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req22_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req22_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req22_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req22_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req22_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req22_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req22_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req22_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req22_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req22_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req22_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req22_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req22_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[23]) begin
		gnt_pre[23] = (req23_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req23_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req23_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req23_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req23_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req23_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req23_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req23_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req23_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req23_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req23_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req23_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req23_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req23_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req23_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req23_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req23_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req23_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req23_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req23_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req23_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req23_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req23_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req23_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req23_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req23_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req23_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req23_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req23_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req23_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req23_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req23_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req23_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req23_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req23_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req23_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req23_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req23_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req23_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req23_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req23_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req23_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req23_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req23_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req23_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req23_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req23_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req23_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req23_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req23_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req23_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req23_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req23_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req23_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req23_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req23_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req23_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req23_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req23_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req23_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req23_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req23_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req23_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req23_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[24]) begin
		gnt_pre[24] = (req24_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req24_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req24_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req24_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req24_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req24_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req24_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req24_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req24_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req24_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req24_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req24_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req24_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req24_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req24_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req24_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req24_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req24_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req24_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req24_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req24_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req24_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req24_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req24_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req24_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req24_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req24_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req24_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req24_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req24_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req24_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req24_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req24_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req24_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req24_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req24_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req24_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req24_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req24_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req24_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req24_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req24_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req24_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req24_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req24_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req24_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req24_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req24_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req24_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req24_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req24_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req24_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req24_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req24_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req24_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req24_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req24_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req24_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req24_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req24_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req24_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req24_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req24_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req24_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[25]) begin
		gnt_pre[25] = (req25_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req25_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req25_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req25_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req25_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req25_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req25_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req25_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req25_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req25_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req25_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req25_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req25_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req25_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req25_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req25_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req25_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req25_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req25_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req25_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req25_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req25_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req25_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req25_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req25_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req25_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req25_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req25_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req25_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req25_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req25_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req25_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req25_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req25_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req25_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req25_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req25_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req25_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req25_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req25_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req25_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req25_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req25_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req25_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req25_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req25_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req25_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req25_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req25_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req25_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req25_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req25_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req25_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req25_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req25_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req25_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req25_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req25_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req25_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req25_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req25_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req25_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req25_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req25_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[26]) begin
		gnt_pre[26] = (req26_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req26_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req26_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req26_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req26_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req26_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req26_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req26_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req26_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req26_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req26_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req26_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req26_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req26_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req26_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req26_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req26_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req26_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req26_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req26_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req26_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req26_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req26_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req26_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req26_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req26_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req26_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req26_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req26_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req26_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req26_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req26_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req26_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req26_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req26_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req26_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req26_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req26_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req26_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req26_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req26_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req26_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req26_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req26_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req26_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req26_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req26_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req26_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req26_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req26_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req26_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req26_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req26_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req26_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req26_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req26_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req26_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req26_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req26_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req26_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req26_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req26_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req26_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req26_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[27]) begin
		gnt_pre[27] = (req27_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req27_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req27_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req27_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req27_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req27_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req27_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req27_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req27_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req27_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req27_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req27_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req27_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req27_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req27_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req27_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req27_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req27_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req27_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req27_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req27_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req27_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req27_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req27_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req27_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req27_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req27_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req27_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req27_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req27_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req27_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req27_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req27_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req27_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req27_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req27_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req27_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req27_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req27_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req27_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req27_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req27_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req27_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req27_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req27_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req27_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req27_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req27_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req27_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req27_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req27_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req27_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req27_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req27_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req27_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req27_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req27_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req27_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req27_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req27_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req27_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req27_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req27_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req27_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[28]) begin
		gnt_pre[28] = (req28_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req28_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req28_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req28_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req28_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req28_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req28_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req28_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req28_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req28_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req28_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req28_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req28_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req28_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req28_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req28_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req28_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req28_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req28_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req28_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req28_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req28_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req28_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req28_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req28_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req28_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req28_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req28_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req28_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req28_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req28_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req28_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req28_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req28_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req28_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req28_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req28_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req28_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req28_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req28_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req28_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req28_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req28_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req28_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req28_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req28_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req28_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req28_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req28_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req28_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req28_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req28_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req28_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req28_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req28_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req28_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req28_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req28_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req28_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req28_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req28_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req28_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req28_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req28_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[29]) begin
		gnt_pre[29] = (req29_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req29_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req29_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req29_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req29_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req29_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req29_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req29_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req29_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req29_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req29_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req29_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req29_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req29_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req29_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req29_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req29_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req29_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req29_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req29_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req29_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req29_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req29_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req29_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req29_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req29_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req29_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req29_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req29_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req29_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req29_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req29_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req29_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req29_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req29_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req29_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req29_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req29_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req29_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req29_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req29_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req29_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req29_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req29_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req29_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req29_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req29_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req29_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req29_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req29_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req29_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req29_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req29_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req29_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req29_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req29_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req29_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req29_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req29_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req29_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req29_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req29_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req29_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req29_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[30]) begin
		gnt_pre[30] = (req30_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req30_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req30_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req30_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req30_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req30_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req30_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req30_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req30_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req30_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req30_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req30_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req30_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req30_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req30_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req30_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req30_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req30_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req30_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req30_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req30_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req30_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req30_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req30_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req30_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req30_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req30_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req30_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req30_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req30_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req30_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req30_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req30_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req30_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req30_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req30_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req30_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req30_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req30_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req30_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req30_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req30_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req30_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req30_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req30_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req30_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req30_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req30_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req30_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req30_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req30_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req30_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req30_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req30_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req30_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req30_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req30_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req30_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req30_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req30_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req30_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req30_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req30_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req30_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[31]) begin
		gnt_pre[31] = (req31_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req31_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req31_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req31_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req31_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req31_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req31_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req31_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req31_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req31_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req31_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req31_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req31_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req31_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req31_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req31_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req31_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req31_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req31_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req31_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req31_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req31_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req31_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req31_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req31_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req31_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req31_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req31_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req31_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req31_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req31_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req31_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req31_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req31_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req31_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req31_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req31_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req31_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req31_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req31_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req31_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req31_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req31_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req31_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req31_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req31_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req31_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req31_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req31_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req31_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req31_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req31_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req31_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req31_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req31_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req31_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req31_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req31_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req31_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req31_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req31_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req31_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req31_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req31_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[32]) begin
		gnt_pre[32] = (req32_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req32_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req32_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req32_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req32_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req32_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req32_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req32_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req32_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req32_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req32_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req32_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req32_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req32_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req32_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req32_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req32_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req32_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req32_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req32_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req32_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req32_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req32_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req32_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req32_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req32_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req32_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req32_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req32_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req32_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req32_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req32_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req32_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req32_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req32_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req32_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req32_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req32_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req32_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req32_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req32_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req32_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req32_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req32_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req32_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req32_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req32_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req32_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req32_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req32_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req32_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req32_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req32_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req32_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req32_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req32_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req32_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req32_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req32_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req32_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req32_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req32_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req32_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req32_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[33]) begin
		gnt_pre[33] = (req33_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req33_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req33_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req33_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req33_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req33_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req33_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req33_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req33_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req33_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req33_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req33_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req33_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req33_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req33_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req33_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req33_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req33_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req33_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req33_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req33_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req33_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req33_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req33_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req33_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req33_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req33_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req33_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req33_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req33_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req33_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req33_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req33_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req33_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req33_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req33_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req33_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req33_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req33_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req33_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req33_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req33_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req33_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req33_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req33_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req33_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req33_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req33_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req33_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req33_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req33_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req33_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req33_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req33_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req33_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req33_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req33_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req33_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req33_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req33_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req33_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req33_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req33_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req33_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[34]) begin
		gnt_pre[34] = (req34_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req34_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req34_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req34_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req34_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req34_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req34_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req34_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req34_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req34_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req34_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req34_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req34_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req34_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req34_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req34_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req34_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req34_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req34_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req34_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req34_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req34_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req34_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req34_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req34_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req34_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req34_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req34_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req34_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req34_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req34_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req34_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req34_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req34_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req34_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req34_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req34_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req34_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req34_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req34_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req34_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req34_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req34_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req34_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req34_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req34_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req34_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req34_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req34_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req34_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req34_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req34_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req34_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req34_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req34_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req34_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req34_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req34_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req34_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req34_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req34_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req34_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req34_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req34_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[35]) begin
		gnt_pre[35] = (req35_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req35_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req35_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req35_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req35_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req35_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req35_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req35_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req35_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req35_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req35_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req35_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req35_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req35_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req35_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req35_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req35_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req35_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req35_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req35_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req35_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req35_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req35_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req35_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req35_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req35_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req35_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req35_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req35_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req35_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req35_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req35_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req35_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req35_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req35_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req35_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req35_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req35_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req35_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req35_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req35_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req35_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req35_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req35_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req35_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req35_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req35_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req35_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req35_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req35_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req35_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req35_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req35_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req35_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req35_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req35_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req35_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req35_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req35_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req35_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req35_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req35_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req35_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req35_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[36]) begin
		gnt_pre[36] = (req36_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req36_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req36_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req36_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req36_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req36_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req36_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req36_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req36_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req36_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req36_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req36_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req36_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req36_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req36_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req36_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req36_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req36_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req36_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req36_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req36_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req36_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req36_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req36_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req36_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req36_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req36_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req36_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req36_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req36_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req36_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req36_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req36_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req36_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req36_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req36_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req36_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req36_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req36_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req36_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req36_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req36_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req36_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req36_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req36_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req36_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req36_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req36_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req36_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req36_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req36_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req36_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req36_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req36_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req36_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req36_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req36_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req36_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req36_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req36_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req36_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req36_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req36_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req36_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[37]) begin
		gnt_pre[37] = (req37_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req37_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req37_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req37_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req37_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req37_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req37_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req37_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req37_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req37_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req37_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req37_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req37_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req37_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req37_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req37_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req37_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req37_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req37_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req37_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req37_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req37_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req37_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req37_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req37_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req37_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req37_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req37_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req37_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req37_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req37_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req37_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req37_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req37_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req37_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req37_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req37_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req37_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req37_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req37_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req37_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req37_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req37_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req37_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req37_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req37_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req37_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req37_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req37_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req37_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req37_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req37_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req37_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req37_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req37_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req37_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req37_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req37_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req37_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req37_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req37_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req37_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req37_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req37_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[38]) begin
		gnt_pre[38] = (req38_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req38_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req38_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req38_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req38_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req38_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req38_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req38_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req38_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req38_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req38_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req38_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req38_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req38_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req38_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req38_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req38_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req38_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req38_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req38_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req38_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req38_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req38_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req38_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req38_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req38_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req38_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req38_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req38_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req38_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req38_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req38_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req38_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req38_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req38_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req38_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req38_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req38_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req38_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req38_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req38_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req38_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req38_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req38_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req38_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req38_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req38_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req38_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req38_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req38_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req38_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req38_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req38_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req38_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req38_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req38_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req38_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req38_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req38_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req38_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req38_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req38_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req38_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req38_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[39]) begin
		gnt_pre[39] = (req39_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req39_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req39_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req39_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req39_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req39_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req39_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req39_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req39_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req39_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req39_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req39_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req39_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req39_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req39_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req39_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req39_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req39_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req39_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req39_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req39_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req39_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req39_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req39_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req39_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req39_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req39_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req39_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req39_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req39_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req39_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req39_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req39_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req39_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req39_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req39_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req39_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req39_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req39_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req39_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req39_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req39_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req39_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req39_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req39_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req39_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req39_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req39_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req39_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req39_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req39_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req39_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req39_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req39_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req39_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req39_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req39_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req39_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req39_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req39_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req39_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req39_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req39_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req39_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[40]) begin
		gnt_pre[40] = (req40_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req40_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req40_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req40_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req40_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req40_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req40_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req40_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req40_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req40_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req40_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req40_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req40_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req40_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req40_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req40_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req40_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req40_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req40_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req40_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req40_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req40_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req40_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req40_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req40_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req40_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req40_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req40_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req40_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req40_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req40_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req40_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req40_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req40_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req40_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req40_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req40_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req40_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req40_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req40_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req40_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req40_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req40_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req40_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req40_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req40_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req40_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req40_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req40_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req40_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req40_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req40_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req40_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req40_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req40_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req40_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req40_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req40_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req40_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req40_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req40_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req40_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req40_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req40_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[41]) begin
		gnt_pre[41] = (req41_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req41_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req41_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req41_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req41_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req41_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req41_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req41_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req41_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req41_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req41_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req41_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req41_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req41_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req41_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req41_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req41_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req41_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req41_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req41_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req41_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req41_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req41_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req41_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req41_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req41_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req41_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req41_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req41_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req41_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req41_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req41_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req41_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req41_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req41_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req41_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req41_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req41_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req41_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req41_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req41_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req41_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req41_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req41_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req41_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req41_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req41_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req41_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req41_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req41_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req41_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req41_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req41_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req41_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req41_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req41_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req41_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req41_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req41_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req41_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req41_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req41_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req41_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req41_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[42]) begin
		gnt_pre[42] = (req42_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req42_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req42_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req42_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req42_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req42_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req42_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req42_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req42_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req42_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req42_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req42_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req42_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req42_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req42_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req42_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req42_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req42_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req42_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req42_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req42_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req42_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req42_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req42_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req42_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req42_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req42_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req42_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req42_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req42_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req42_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req42_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req42_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req42_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req42_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req42_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req42_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req42_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req42_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req42_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req42_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req42_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req42_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req42_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req42_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req42_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req42_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req42_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req42_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req42_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req42_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req42_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req42_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req42_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req42_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req42_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req42_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req42_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req42_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req42_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req42_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req42_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req42_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req42_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[43]) begin
		gnt_pre[43] = (req43_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req43_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req43_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req43_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req43_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req43_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req43_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req43_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req43_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req43_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req43_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req43_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req43_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req43_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req43_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req43_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req43_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req43_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req43_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req43_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req43_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req43_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req43_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req43_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req43_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req43_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req43_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req43_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req43_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req43_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req43_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req43_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req43_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req43_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req43_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req43_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req43_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req43_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req43_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req43_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req43_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req43_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req43_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req43_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req43_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req43_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req43_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req43_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req43_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req43_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req43_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req43_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req43_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req43_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req43_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req43_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req43_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req43_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req43_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req43_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req43_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req43_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req43_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req43_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[44]) begin
		gnt_pre[44] = (req44_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req44_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req44_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req44_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req44_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req44_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req44_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req44_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req44_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req44_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req44_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req44_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req44_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req44_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req44_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req44_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req44_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req44_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req44_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req44_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req44_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req44_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req44_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req44_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req44_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req44_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req44_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req44_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req44_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req44_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req44_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req44_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req44_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req44_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req44_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req44_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req44_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req44_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req44_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req44_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req44_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req44_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req44_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req44_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req44_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req44_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req44_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req44_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req44_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req44_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req44_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req44_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req44_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req44_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req44_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req44_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req44_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req44_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req44_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req44_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req44_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req44_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req44_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req44_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[45]) begin
		gnt_pre[45] = (req45_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req45_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req45_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req45_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req45_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req45_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req45_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req45_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req45_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req45_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req45_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req45_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req45_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req45_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req45_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req45_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req45_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req45_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req45_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req45_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req45_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req45_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req45_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req45_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req45_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req45_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req45_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req45_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req45_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req45_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req45_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req45_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req45_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req45_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req45_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req45_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req45_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req45_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req45_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req45_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req45_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req45_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req45_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req45_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req45_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req45_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req45_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req45_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req45_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req45_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req45_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req45_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req45_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req45_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req45_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req45_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req45_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req45_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req45_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req45_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req45_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req45_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req45_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req45_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[46]) begin
		gnt_pre[46] = (req46_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req46_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req46_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req46_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req46_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req46_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req46_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req46_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req46_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req46_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req46_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req46_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req46_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req46_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req46_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req46_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req46_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req46_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req46_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req46_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req46_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req46_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req46_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req46_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req46_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req46_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req46_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req46_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req46_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req46_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req46_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req46_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req46_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req46_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req46_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req46_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req46_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req46_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req46_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req46_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req46_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req46_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req46_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req46_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req46_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req46_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req46_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req46_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req46_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req46_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req46_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req46_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req46_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req46_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req46_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req46_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req46_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req46_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req46_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req46_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req46_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req46_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req46_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req46_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[47]) begin
		gnt_pre[47] = (req47_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req47_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req47_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req47_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req47_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req47_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req47_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req47_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req47_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req47_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req47_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req47_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req47_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req47_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req47_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req47_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req47_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req47_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req47_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req47_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req47_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req47_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req47_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req47_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req47_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req47_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req47_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req47_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req47_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req47_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req47_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req47_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req47_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req47_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req47_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req47_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req47_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req47_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req47_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req47_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req47_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req47_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req47_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req47_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req47_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req47_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req47_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req47_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req47_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req47_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req47_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req47_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req47_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req47_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req47_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req47_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req47_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req47_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req47_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req47_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req47_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req47_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req47_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req47_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[48]) begin
		gnt_pre[48] = (req48_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req48_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req48_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req48_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req48_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req48_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req48_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req48_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req48_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req48_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req48_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req48_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req48_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req48_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req48_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req48_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req48_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req48_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req48_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req48_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req48_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req48_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req48_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req48_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req48_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req48_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req48_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req48_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req48_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req48_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req48_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req48_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req48_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req48_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req48_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req48_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req48_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req48_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req48_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req48_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req48_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req48_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req48_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req48_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req48_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req48_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req48_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req48_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req48_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req48_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req48_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req48_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req48_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req48_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req48_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req48_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req48_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req48_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req48_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req48_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req48_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req48_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req48_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req48_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[49]) begin
		gnt_pre[49] = (req49_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req49_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req49_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req49_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req49_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req49_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req49_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req49_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req49_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req49_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req49_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req49_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req49_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req49_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req49_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req49_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req49_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req49_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req49_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req49_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req49_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req49_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req49_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req49_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req49_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req49_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req49_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req49_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req49_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req49_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req49_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req49_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req49_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req49_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req49_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req49_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req49_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req49_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req49_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req49_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req49_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req49_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req49_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req49_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req49_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req49_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req49_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req49_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req49_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req49_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req49_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req49_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req49_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req49_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req49_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req49_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req49_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req49_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req49_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req49_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req49_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req49_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req49_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req49_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[50]) begin
		gnt_pre[50] = (req50_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req50_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req50_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req50_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req50_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req50_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req50_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req50_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req50_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req50_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req50_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req50_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req50_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req50_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req50_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req50_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req50_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req50_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req50_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req50_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req50_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req50_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req50_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req50_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req50_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req50_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req50_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req50_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req50_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req50_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req50_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req50_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req50_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req50_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req50_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req50_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req50_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req50_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req50_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req50_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req50_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req50_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req50_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req50_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req50_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req50_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req50_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req50_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req50_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req50_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req50_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req50_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req50_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req50_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req50_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req50_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req50_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req50_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req50_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req50_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req50_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req50_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req50_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req50_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[51]) begin
		gnt_pre[51] = (req51_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req51_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req51_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req51_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req51_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req51_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req51_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req51_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req51_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req51_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req51_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req51_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req51_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req51_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req51_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req51_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req51_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req51_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req51_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req51_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req51_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req51_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req51_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req51_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req51_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req51_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req51_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req51_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req51_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req51_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req51_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req51_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req51_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req51_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req51_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req51_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req51_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req51_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req51_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req51_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req51_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req51_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req51_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req51_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req51_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req51_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req51_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req51_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req51_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req51_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req51_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req51_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req51_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req51_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req51_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req51_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req51_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req51_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req51_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req51_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req51_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req51_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req51_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req51_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[52]) begin
		gnt_pre[52] = (req52_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req52_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req52_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req52_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req52_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req52_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req52_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req52_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req52_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req52_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req52_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req52_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req52_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req52_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req52_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req52_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req52_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req52_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req52_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req52_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req52_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req52_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req52_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req52_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req52_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req52_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req52_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req52_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req52_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req52_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req52_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req52_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req52_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req52_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req52_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req52_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req52_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req52_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req52_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req52_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req52_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req52_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req52_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req52_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req52_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req52_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req52_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req52_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req52_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req52_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req52_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req52_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req52_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req52_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req52_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req52_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req52_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req52_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req52_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req52_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req52_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req52_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req52_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req52_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[53]) begin
		gnt_pre[53] = (req53_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req53_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req53_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req53_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req53_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req53_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req53_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req53_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req53_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req53_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req53_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req53_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req53_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req53_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req53_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req53_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req53_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req53_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req53_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req53_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req53_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req53_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req53_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req53_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req53_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req53_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req53_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req53_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req53_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req53_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req53_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req53_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req53_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req53_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req53_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req53_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req53_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req53_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req53_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req53_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req53_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req53_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req53_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req53_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req53_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req53_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req53_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req53_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req53_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req53_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req53_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req53_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req53_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req53_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req53_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req53_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req53_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req53_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req53_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req53_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req53_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req53_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req53_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req53_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[54]) begin
		gnt_pre[54] = (req54_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req54_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req54_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req54_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req54_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req54_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req54_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req54_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req54_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req54_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req54_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req54_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req54_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req54_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req54_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req54_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req54_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req54_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req54_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req54_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req54_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req54_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req54_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req54_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req54_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req54_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req54_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req54_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req54_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req54_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req54_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req54_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req54_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req54_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req54_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req54_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req54_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req54_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req54_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req54_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req54_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req54_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req54_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req54_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req54_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req54_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req54_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req54_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req54_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req54_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req54_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req54_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req54_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req54_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req54_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req54_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req54_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req54_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req54_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req54_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req54_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req54_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req54_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req54_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[55]) begin
		gnt_pre[55] = (req55_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req55_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req55_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req55_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req55_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req55_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req55_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req55_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req55_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req55_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req55_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req55_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req55_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req55_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req55_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req55_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req55_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req55_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req55_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req55_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req55_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req55_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req55_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req55_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req55_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req55_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req55_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req55_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req55_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req55_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req55_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req55_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req55_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req55_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req55_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req55_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req55_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req55_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req55_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req55_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req55_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req55_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req55_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req55_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req55_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req55_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req55_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req55_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req55_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req55_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req55_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req55_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req55_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req55_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req55_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req55_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req55_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req55_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req55_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req55_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req55_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req55_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req55_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req55_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[56]) begin
		gnt_pre[56] = (req56_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req56_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req56_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req56_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req56_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req56_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req56_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req56_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req56_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req56_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req56_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req56_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req56_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req56_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req56_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req56_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req56_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req56_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req56_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req56_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req56_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req56_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req56_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req56_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req56_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req56_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req56_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req56_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req56_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req56_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req56_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req56_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req56_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req56_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req56_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req56_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req56_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req56_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req56_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req56_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req56_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req56_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req56_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req56_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req56_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req56_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req56_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req56_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req56_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req56_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req56_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req56_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req56_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req56_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req56_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req56_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req56_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req56_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req56_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req56_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req56_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req56_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req56_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req56_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[57]) begin
		gnt_pre[57] = (req57_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req57_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req57_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req57_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req57_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req57_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req57_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req57_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req57_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req57_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req57_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req57_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req57_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req57_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req57_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req57_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req57_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req57_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req57_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req57_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req57_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req57_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req57_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req57_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req57_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req57_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req57_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req57_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req57_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req57_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req57_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req57_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req57_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req57_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req57_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req57_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req57_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req57_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req57_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req57_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req57_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req57_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req57_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req57_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req57_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req57_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req57_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req57_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req57_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req57_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req57_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req57_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req57_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req57_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req57_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req57_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req57_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req57_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req57_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req57_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req57_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req57_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req57_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req57_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[58]) begin
		gnt_pre[58] = (req58_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req58_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req58_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req58_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req58_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req58_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req58_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req58_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req58_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req58_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req58_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req58_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req58_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req58_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req58_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req58_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req58_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req58_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req58_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req58_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req58_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req58_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req58_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req58_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req58_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req58_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req58_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req58_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req58_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req58_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req58_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req58_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req58_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req58_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req58_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req58_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req58_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req58_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req58_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req58_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req58_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req58_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req58_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req58_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req58_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req58_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req58_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req58_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req58_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req58_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req58_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req58_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req58_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req58_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req58_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req58_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req58_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req58_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req58_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req58_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req58_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req58_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req58_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req58_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[59]) begin
		gnt_pre[59] = (req59_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req59_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req59_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req59_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req59_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req59_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req59_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req59_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req59_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req59_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req59_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req59_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req59_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req59_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req59_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req59_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req59_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req59_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req59_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req59_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req59_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req59_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req59_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req59_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req59_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req59_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req59_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req59_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req59_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req59_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req59_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req59_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req59_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req59_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req59_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req59_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req59_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req59_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req59_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req59_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req59_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req59_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req59_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req59_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req59_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req59_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req59_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req59_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req59_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req59_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req59_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req59_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req59_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req59_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req59_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req59_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req59_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req59_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req59_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req59_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req59_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req59_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req59_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req59_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[60]) begin
		gnt_pre[60] = (req60_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req60_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req60_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req60_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req60_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req60_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req60_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req60_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req60_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req60_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req60_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req60_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req60_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req60_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req60_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req60_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req60_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req60_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req60_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req60_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req60_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req60_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req60_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req60_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req60_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req60_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req60_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req60_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req60_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req60_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req60_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req60_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req60_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req60_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req60_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req60_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req60_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req60_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req60_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req60_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req60_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req60_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req60_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req60_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req60_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req60_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req60_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req60_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req60_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req60_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req60_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req60_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req60_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req60_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req60_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req60_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req60_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req60_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req60_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req60_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req60_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req60_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req60_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req60_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[61]) begin
		gnt_pre[61] = (req61_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req61_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req61_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req61_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req61_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req61_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req61_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req61_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req61_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req61_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req61_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req61_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req61_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req61_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req61_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req61_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req61_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req61_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req61_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req61_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req61_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req61_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req61_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req61_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req61_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req61_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req61_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req61_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req61_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req61_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req61_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req61_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req61_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req61_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req61_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req61_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req61_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req61_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req61_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req61_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req61_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req61_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req61_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req61_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req61_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req61_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req61_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req61_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req61_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req61_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req61_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req61_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req61_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req61_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req61_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req61_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req61_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req61_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req61_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req61_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req61_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req61_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req61_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req61_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[62]) begin
		gnt_pre[62] = (req62_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req62_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req62_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req62_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req62_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req62_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req62_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req62_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req62_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req62_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req62_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req62_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req62_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req62_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req62_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req62_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req62_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req62_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req62_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req62_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req62_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req62_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req62_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req62_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req62_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req62_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req62_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req62_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req62_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req62_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req62_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req62_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req62_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req62_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req62_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req62_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req62_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req62_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req62_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req62_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req62_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req62_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req62_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req62_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req62_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req62_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req62_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req62_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req62_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req62_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req62_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req62_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req62_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req62_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req62_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req62_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req62_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req62_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req62_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req62_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req62_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req62_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req62_used_status)) ?1'b0 |
	((req63 & (req63_used_status > req62_used_status)) ?1'b0 |
		1'b1;
	end
	if(req[63]) begin
		gnt_pre[63] = (req63_used_status==64) ? 1'b1 |

	((req0 & (req0_used_status > req63_used_status)) ?1'b0 |
	((req1 & (req1_used_status > req63_used_status)) ?1'b0 |
	((req2 & (req2_used_status > req63_used_status)) ?1'b0 |
	((req3 & (req3_used_status > req63_used_status)) ?1'b0 |
	((req4 & (req4_used_status > req63_used_status)) ?1'b0 |
	((req5 & (req5_used_status > req63_used_status)) ?1'b0 |
	((req6 & (req6_used_status > req63_used_status)) ?1'b0 |
	((req7 & (req7_used_status > req63_used_status)) ?1'b0 |
	((req8 & (req8_used_status > req63_used_status)) ?1'b0 |
	((req9 & (req9_used_status > req63_used_status)) ?1'b0 |
	((req10 & (req10_used_status > req63_used_status)) ?1'b0 |
	((req11 & (req11_used_status > req63_used_status)) ?1'b0 |
	((req12 & (req12_used_status > req63_used_status)) ?1'b0 |
	((req13 & (req13_used_status > req63_used_status)) ?1'b0 |
	((req14 & (req14_used_status > req63_used_status)) ?1'b0 |
	((req15 & (req15_used_status > req63_used_status)) ?1'b0 |
	((req16 & (req16_used_status > req63_used_status)) ?1'b0 |
	((req17 & (req17_used_status > req63_used_status)) ?1'b0 |
	((req18 & (req18_used_status > req63_used_status)) ?1'b0 |
	((req19 & (req19_used_status > req63_used_status)) ?1'b0 |
	((req20 & (req20_used_status > req63_used_status)) ?1'b0 |
	((req21 & (req21_used_status > req63_used_status)) ?1'b0 |
	((req22 & (req22_used_status > req63_used_status)) ?1'b0 |
	((req23 & (req23_used_status > req63_used_status)) ?1'b0 |
	((req24 & (req24_used_status > req63_used_status)) ?1'b0 |
	((req25 & (req25_used_status > req63_used_status)) ?1'b0 |
	((req26 & (req26_used_status > req63_used_status)) ?1'b0 |
	((req27 & (req27_used_status > req63_used_status)) ?1'b0 |
	((req28 & (req28_used_status > req63_used_status)) ?1'b0 |
	((req29 & (req29_used_status > req63_used_status)) ?1'b0 |
	((req30 & (req30_used_status > req63_used_status)) ?1'b0 |
	((req31 & (req31_used_status > req63_used_status)) ?1'b0 |
	((req32 & (req32_used_status > req63_used_status)) ?1'b0 |
	((req33 & (req33_used_status > req63_used_status)) ?1'b0 |
	((req34 & (req34_used_status > req63_used_status)) ?1'b0 |
	((req35 & (req35_used_status > req63_used_status)) ?1'b0 |
	((req36 & (req36_used_status > req63_used_status)) ?1'b0 |
	((req37 & (req37_used_status > req63_used_status)) ?1'b0 |
	((req38 & (req38_used_status > req63_used_status)) ?1'b0 |
	((req39 & (req39_used_status > req63_used_status)) ?1'b0 |
	((req40 & (req40_used_status > req63_used_status)) ?1'b0 |
	((req41 & (req41_used_status > req63_used_status)) ?1'b0 |
	((req42 & (req42_used_status > req63_used_status)) ?1'b0 |
	((req43 & (req43_used_status > req63_used_status)) ?1'b0 |
	((req44 & (req44_used_status > req63_used_status)) ?1'b0 |
	((req45 & (req45_used_status > req63_used_status)) ?1'b0 |
	((req46 & (req46_used_status > req63_used_status)) ?1'b0 |
	((req47 & (req47_used_status > req63_used_status)) ?1'b0 |
	((req48 & (req48_used_status > req63_used_status)) ?1'b0 |
	((req49 & (req49_used_status > req63_used_status)) ?1'b0 |
	((req50 & (req50_used_status > req63_used_status)) ?1'b0 |
	((req51 & (req51_used_status > req63_used_status)) ?1'b0 |
	((req52 & (req52_used_status > req63_used_status)) ?1'b0 |
	((req53 & (req53_used_status > req63_used_status)) ?1'b0 |
	((req54 & (req54_used_status > req63_used_status)) ?1'b0 |
	((req55 & (req55_used_status > req63_used_status)) ?1'b0 |
	((req56 & (req56_used_status > req63_used_status)) ?1'b0 |
	((req57 & (req57_used_status > req63_used_status)) ?1'b0 |
	((req58 & (req58_used_status > req63_used_status)) ?1'b0 |
	((req59 & (req59_used_status > req63_used_status)) ?1'b0 |
	((req60 & (req60_used_status > req63_used_status)) ?1'b0 |
	((req61 & (req61_used_status > req63_used_status)) ?1'b0 |
	((req62 & (req62_used_status > req63_used_status)) ?1'b0 |
		1'b1;
	end

assign gnt[63:0] = gnt_pre[63:0];

endmodule
