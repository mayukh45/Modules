
module AH_demux_12_258_0 (select
,ing_data
,ing_valid
,ing_ready
,egr0_data
,egr0_valid
,egr0_ready
,egr1_data
,egr1_valid
,egr1_ready
,egr2_data
,egr2_valid
,egr2_ready
,egr3_data
,egr3_valid
,egr3_ready
,egr4_data
,egr4_valid
,egr4_ready
,egr5_data
,egr5_valid
,egr5_ready
,egr6_data
,egr6_valid
,egr6_ready
,egr7_data
,egr7_valid
,egr7_ready
,egr8_data
,egr8_valid
,egr8_ready
,egr9_data
,egr9_valid
,egr9_ready
,egr10_data
,egr10_valid
,egr10_ready
,egr11_data
,egr11_valid
,egr11_ready
,egr12_data
,egr12_valid
,egr12_ready
,egr13_data
,egr13_valid
,egr13_ready
,egr14_data
,egr14_valid
,egr14_ready
,egr15_data
,egr15_valid
,egr15_ready
,egr16_data
,egr16_valid
,egr16_ready
,egr17_data
,egr17_valid
,egr17_ready
,egr18_data
,egr18_valid
,egr18_ready
,egr19_data
,egr19_valid
,egr19_ready
,egr20_data
,egr20_valid
,egr20_ready
,egr21_data
,egr21_valid
,egr21_ready
,egr22_data
,egr22_valid
,egr22_ready
,egr23_data
,egr23_valid
,egr23_ready
,egr24_data
,egr24_valid
,egr24_ready
,egr25_data
,egr25_valid
,egr25_ready
,egr26_data
,egr26_valid
,egr26_ready
,egr27_data
,egr27_valid
,egr27_ready
,egr28_data
,egr28_valid
,egr28_ready
,egr29_data
,egr29_valid
,egr29_ready
,egr30_data
,egr30_valid
,egr30_ready
,egr31_data
,egr31_valid
,egr31_ready
,egr32_data
,egr32_valid
,egr32_ready
,egr33_data
,egr33_valid
,egr33_ready
,egr34_data
,egr34_valid
,egr34_ready
,egr35_data
,egr35_valid
,egr35_ready
,egr36_data
,egr36_valid
,egr36_ready
,egr37_data
,egr37_valid
,egr37_ready
,egr38_data
,egr38_valid
,egr38_ready
,egr39_data
,egr39_valid
,egr39_ready
,egr40_data
,egr40_valid
,egr40_ready
,egr41_data
,egr41_valid
,egr41_ready
,egr42_data
,egr42_valid
,egr42_ready
,egr43_data
,egr43_valid
,egr43_ready
,egr44_data
,egr44_valid
,egr44_ready
,egr45_data
,egr45_valid
,egr45_ready
,egr46_data
,egr46_valid
,egr46_ready
,egr47_data
,egr47_valid
,egr47_ready
,egr48_data
,egr48_valid
,egr48_ready
,egr49_data
,egr49_valid
,egr49_ready
,egr50_data
,egr50_valid
,egr50_ready
,egr51_data
,egr51_valid
,egr51_ready
,egr52_data
,egr52_valid
,egr52_ready
,egr53_data
,egr53_valid
,egr53_ready
,egr54_data
,egr54_valid
,egr54_ready
,egr55_data
,egr55_valid
,egr55_ready
,egr56_data
,egr56_valid
,egr56_ready
,egr57_data
,egr57_valid
,egr57_ready
,egr58_data
,egr58_valid
,egr58_ready
,egr59_data
,egr59_valid
,egr59_ready
,egr60_data
,egr60_valid
,egr60_ready
,egr61_data
,egr61_valid
,egr61_ready
,egr62_data
,egr62_valid
,egr62_ready
,egr63_data
,egr63_valid
,egr63_ready
,egr64_data
,egr64_valid
,egr64_ready
,egr65_data
,egr65_valid
,egr65_ready
,egr66_data
,egr66_valid
,egr66_ready
,egr67_data
,egr67_valid
,egr67_ready
,egr68_data
,egr68_valid
,egr68_ready
,egr69_data
,egr69_valid
,egr69_ready
,egr70_data
,egr70_valid
,egr70_ready
,egr71_data
,egr71_valid
,egr71_ready
,egr72_data
,egr72_valid
,egr72_ready
,egr73_data
,egr73_valid
,egr73_ready
,egr74_data
,egr74_valid
,egr74_ready
,egr75_data
,egr75_valid
,egr75_ready
,egr76_data
,egr76_valid
,egr76_ready
,egr77_data
,egr77_valid
,egr77_ready
,egr78_data
,egr78_valid
,egr78_ready
,egr79_data
,egr79_valid
,egr79_ready
,egr80_data
,egr80_valid
,egr80_ready
,egr81_data
,egr81_valid
,egr81_ready
,egr82_data
,egr82_valid
,egr82_ready
,egr83_data
,egr83_valid
,egr83_ready
,egr84_data
,egr84_valid
,egr84_ready
,egr85_data
,egr85_valid
,egr85_ready
,egr86_data
,egr86_valid
,egr86_ready
,egr87_data
,egr87_valid
,egr87_ready
,egr88_data
,egr88_valid
,egr88_ready
,egr89_data
,egr89_valid
,egr89_ready
,egr90_data
,egr90_valid
,egr90_ready
,egr91_data
,egr91_valid
,egr91_ready
,egr92_data
,egr92_valid
,egr92_ready
,egr93_data
,egr93_valid
,egr93_ready
,egr94_data
,egr94_valid
,egr94_ready
,egr95_data
,egr95_valid
,egr95_ready
,egr96_data
,egr96_valid
,egr96_ready
,egr97_data
,egr97_valid
,egr97_ready
,egr98_data
,egr98_valid
,egr98_ready
,egr99_data
,egr99_valid
,egr99_ready
,egr100_data
,egr100_valid
,egr100_ready
,egr101_data
,egr101_valid
,egr101_ready
,egr102_data
,egr102_valid
,egr102_ready
,egr103_data
,egr103_valid
,egr103_ready
,egr104_data
,egr104_valid
,egr104_ready
,egr105_data
,egr105_valid
,egr105_ready
,egr106_data
,egr106_valid
,egr106_ready
,egr107_data
,egr107_valid
,egr107_ready
,egr108_data
,egr108_valid
,egr108_ready
,egr109_data
,egr109_valid
,egr109_ready
,egr110_data
,egr110_valid
,egr110_ready
,egr111_data
,egr111_valid
,egr111_ready
,egr112_data
,egr112_valid
,egr112_ready
,egr113_data
,egr113_valid
,egr113_ready
,egr114_data
,egr114_valid
,egr114_ready
,egr115_data
,egr115_valid
,egr115_ready
,egr116_data
,egr116_valid
,egr116_ready
,egr117_data
,egr117_valid
,egr117_ready
,egr118_data
,egr118_valid
,egr118_ready
,egr119_data
,egr119_valid
,egr119_ready
,egr120_data
,egr120_valid
,egr120_ready
,egr121_data
,egr121_valid
,egr121_ready
,egr122_data
,egr122_valid
,egr122_ready
,egr123_data
,egr123_valid
,egr123_ready
,egr124_data
,egr124_valid
,egr124_ready
,egr125_data
,egr125_valid
,egr125_ready
,egr126_data
,egr126_valid
,egr126_ready
,egr127_data
,egr127_valid
,egr127_ready
,egr128_data
,egr128_valid
,egr128_ready
,egr129_data
,egr129_valid
,egr129_ready
,egr130_data
,egr130_valid
,egr130_ready
,egr131_data
,egr131_valid
,egr131_ready
,egr132_data
,egr132_valid
,egr132_ready
,egr133_data
,egr133_valid
,egr133_ready
,egr134_data
,egr134_valid
,egr134_ready
,egr135_data
,egr135_valid
,egr135_ready
,egr136_data
,egr136_valid
,egr136_ready
,egr137_data
,egr137_valid
,egr137_ready
,egr138_data
,egr138_valid
,egr138_ready
,egr139_data
,egr139_valid
,egr139_ready
,egr140_data
,egr140_valid
,egr140_ready
,egr141_data
,egr141_valid
,egr141_ready
,egr142_data
,egr142_valid
,egr142_ready
,egr143_data
,egr143_valid
,egr143_ready
,egr144_data
,egr144_valid
,egr144_ready
,egr145_data
,egr145_valid
,egr145_ready
,egr146_data
,egr146_valid
,egr146_ready
,egr147_data
,egr147_valid
,egr147_ready
,egr148_data
,egr148_valid
,egr148_ready
,egr149_data
,egr149_valid
,egr149_ready
,egr150_data
,egr150_valid
,egr150_ready
,egr151_data
,egr151_valid
,egr151_ready
,egr152_data
,egr152_valid
,egr152_ready
,egr153_data
,egr153_valid
,egr153_ready
,egr154_data
,egr154_valid
,egr154_ready
,egr155_data
,egr155_valid
,egr155_ready
,egr156_data
,egr156_valid
,egr156_ready
,egr157_data
,egr157_valid
,egr157_ready
,egr158_data
,egr158_valid
,egr158_ready
,egr159_data
,egr159_valid
,egr159_ready
,egr160_data
,egr160_valid
,egr160_ready
,egr161_data
,egr161_valid
,egr161_ready
,egr162_data
,egr162_valid
,egr162_ready
,egr163_data
,egr163_valid
,egr163_ready
,egr164_data
,egr164_valid
,egr164_ready
,egr165_data
,egr165_valid
,egr165_ready
,egr166_data
,egr166_valid
,egr166_ready
,egr167_data
,egr167_valid
,egr167_ready
,egr168_data
,egr168_valid
,egr168_ready
,egr169_data
,egr169_valid
,egr169_ready
,egr170_data
,egr170_valid
,egr170_ready
,egr171_data
,egr171_valid
,egr171_ready
,egr172_data
,egr172_valid
,egr172_ready
,egr173_data
,egr173_valid
,egr173_ready
,egr174_data
,egr174_valid
,egr174_ready
,egr175_data
,egr175_valid
,egr175_ready
,egr176_data
,egr176_valid
,egr176_ready
,egr177_data
,egr177_valid
,egr177_ready
,egr178_data
,egr178_valid
,egr178_ready
,egr179_data
,egr179_valid
,egr179_ready
,egr180_data
,egr180_valid
,egr180_ready
,egr181_data
,egr181_valid
,egr181_ready
,egr182_data
,egr182_valid
,egr182_ready
,egr183_data
,egr183_valid
,egr183_ready
,egr184_data
,egr184_valid
,egr184_ready
,egr185_data
,egr185_valid
,egr185_ready
,egr186_data
,egr186_valid
,egr186_ready
,egr187_data
,egr187_valid
,egr187_ready
,egr188_data
,egr188_valid
,egr188_ready
,egr189_data
,egr189_valid
,egr189_ready
,egr190_data
,egr190_valid
,egr190_ready
,egr191_data
,egr191_valid
,egr191_ready
,egr192_data
,egr192_valid
,egr192_ready
,egr193_data
,egr193_valid
,egr193_ready
,egr194_data
,egr194_valid
,egr194_ready
,egr195_data
,egr195_valid
,egr195_ready
,egr196_data
,egr196_valid
,egr196_ready
,egr197_data
,egr197_valid
,egr197_ready
,egr198_data
,egr198_valid
,egr198_ready
,egr199_data
,egr199_valid
,egr199_ready
,egr200_data
,egr200_valid
,egr200_ready
,egr201_data
,egr201_valid
,egr201_ready
,egr202_data
,egr202_valid
,egr202_ready
,egr203_data
,egr203_valid
,egr203_ready
,egr204_data
,egr204_valid
,egr204_ready
,egr205_data
,egr205_valid
,egr205_ready
,egr206_data
,egr206_valid
,egr206_ready
,egr207_data
,egr207_valid
,egr207_ready
,egr208_data
,egr208_valid
,egr208_ready
,egr209_data
,egr209_valid
,egr209_ready
,egr210_data
,egr210_valid
,egr210_ready
,egr211_data
,egr211_valid
,egr211_ready
,egr212_data
,egr212_valid
,egr212_ready
,egr213_data
,egr213_valid
,egr213_ready
,egr214_data
,egr214_valid
,egr214_ready
,egr215_data
,egr215_valid
,egr215_ready
,egr216_data
,egr216_valid
,egr216_ready
,egr217_data
,egr217_valid
,egr217_ready
,egr218_data
,egr218_valid
,egr218_ready
,egr219_data
,egr219_valid
,egr219_ready
,egr220_data
,egr220_valid
,egr220_ready
,egr221_data
,egr221_valid
,egr221_ready
,egr222_data
,egr222_valid
,egr222_ready
,egr223_data
,egr223_valid
,egr223_ready
,egr224_data
,egr224_valid
,egr224_ready
,egr225_data
,egr225_valid
,egr225_ready
,egr226_data
,egr226_valid
,egr226_ready
,egr227_data
,egr227_valid
,egr227_ready
,egr228_data
,egr228_valid
,egr228_ready
,egr229_data
,egr229_valid
,egr229_ready
,egr230_data
,egr230_valid
,egr230_ready
,egr231_data
,egr231_valid
,egr231_ready
,egr232_data
,egr232_valid
,egr232_ready
,egr233_data
,egr233_valid
,egr233_ready
,egr234_data
,egr234_valid
,egr234_ready
,egr235_data
,egr235_valid
,egr235_ready
,egr236_data
,egr236_valid
,egr236_ready
,egr237_data
,egr237_valid
,egr237_ready
,egr238_data
,egr238_valid
,egr238_ready
,egr239_data
,egr239_valid
,egr239_ready
,egr240_data
,egr240_valid
,egr240_ready
,egr241_data
,egr241_valid
,egr241_ready
,egr242_data
,egr242_valid
,egr242_ready
,egr243_data
,egr243_valid
,egr243_ready
,egr244_data
,egr244_valid
,egr244_ready
,egr245_data
,egr245_valid
,egr245_ready
,egr246_data
,egr246_valid
,egr246_ready
,egr247_data
,egr247_valid
,egr247_ready
,egr248_data
,egr248_valid
,egr248_ready
,egr249_data
,egr249_valid
,egr249_ready
,egr250_data
,egr250_valid
,egr250_ready
,egr251_data
,egr251_valid
,egr251_ready
,egr252_data
,egr252_valid
,egr252_ready
,egr253_data
,egr253_valid
,egr253_ready
,egr254_data
,egr254_valid
,egr254_ready
,egr255_data
,egr255_valid
,egr255_ready
,egr256_data
,egr256_valid
,egr256_ready
,egr257_data
,egr257_valid
,egr257_ready);

input select;
input [11:0] ing_data;
input ing_valid;
output ing_ready;
output [11:0] egr0_data;
output egr0_valid;
input egr0_ready;
output [11:0] egr1_data;
output egr1_valid;
input egr1_ready;
output [11:0] egr2_data;
output egr2_valid;
input egr2_ready;
output [11:0] egr3_data;
output egr3_valid;
input egr3_ready;
output [11:0] egr4_data;
output egr4_valid;
input egr4_ready;
output [11:0] egr5_data;
output egr5_valid;
input egr5_ready;
output [11:0] egr6_data;
output egr6_valid;
input egr6_ready;
output [11:0] egr7_data;
output egr7_valid;
input egr7_ready;
output [11:0] egr8_data;
output egr8_valid;
input egr8_ready;
output [11:0] egr9_data;
output egr9_valid;
input egr9_ready;
output [11:0] egr10_data;
output egr10_valid;
input egr10_ready;
output [11:0] egr11_data;
output egr11_valid;
input egr11_ready;
output [11:0] egr12_data;
output egr12_valid;
input egr12_ready;
output [11:0] egr13_data;
output egr13_valid;
input egr13_ready;
output [11:0] egr14_data;
output egr14_valid;
input egr14_ready;
output [11:0] egr15_data;
output egr15_valid;
input egr15_ready;
output [11:0] egr16_data;
output egr16_valid;
input egr16_ready;
output [11:0] egr17_data;
output egr17_valid;
input egr17_ready;
output [11:0] egr18_data;
output egr18_valid;
input egr18_ready;
output [11:0] egr19_data;
output egr19_valid;
input egr19_ready;
output [11:0] egr20_data;
output egr20_valid;
input egr20_ready;
output [11:0] egr21_data;
output egr21_valid;
input egr21_ready;
output [11:0] egr22_data;
output egr22_valid;
input egr22_ready;
output [11:0] egr23_data;
output egr23_valid;
input egr23_ready;
output [11:0] egr24_data;
output egr24_valid;
input egr24_ready;
output [11:0] egr25_data;
output egr25_valid;
input egr25_ready;
output [11:0] egr26_data;
output egr26_valid;
input egr26_ready;
output [11:0] egr27_data;
output egr27_valid;
input egr27_ready;
output [11:0] egr28_data;
output egr28_valid;
input egr28_ready;
output [11:0] egr29_data;
output egr29_valid;
input egr29_ready;
output [11:0] egr30_data;
output egr30_valid;
input egr30_ready;
output [11:0] egr31_data;
output egr31_valid;
input egr31_ready;
output [11:0] egr32_data;
output egr32_valid;
input egr32_ready;
output [11:0] egr33_data;
output egr33_valid;
input egr33_ready;
output [11:0] egr34_data;
output egr34_valid;
input egr34_ready;
output [11:0] egr35_data;
output egr35_valid;
input egr35_ready;
output [11:0] egr36_data;
output egr36_valid;
input egr36_ready;
output [11:0] egr37_data;
output egr37_valid;
input egr37_ready;
output [11:0] egr38_data;
output egr38_valid;
input egr38_ready;
output [11:0] egr39_data;
output egr39_valid;
input egr39_ready;
output [11:0] egr40_data;
output egr40_valid;
input egr40_ready;
output [11:0] egr41_data;
output egr41_valid;
input egr41_ready;
output [11:0] egr42_data;
output egr42_valid;
input egr42_ready;
output [11:0] egr43_data;
output egr43_valid;
input egr43_ready;
output [11:0] egr44_data;
output egr44_valid;
input egr44_ready;
output [11:0] egr45_data;
output egr45_valid;
input egr45_ready;
output [11:0] egr46_data;
output egr46_valid;
input egr46_ready;
output [11:0] egr47_data;
output egr47_valid;
input egr47_ready;
output [11:0] egr48_data;
output egr48_valid;
input egr48_ready;
output [11:0] egr49_data;
output egr49_valid;
input egr49_ready;
output [11:0] egr50_data;
output egr50_valid;
input egr50_ready;
output [11:0] egr51_data;
output egr51_valid;
input egr51_ready;
output [11:0] egr52_data;
output egr52_valid;
input egr52_ready;
output [11:0] egr53_data;
output egr53_valid;
input egr53_ready;
output [11:0] egr54_data;
output egr54_valid;
input egr54_ready;
output [11:0] egr55_data;
output egr55_valid;
input egr55_ready;
output [11:0] egr56_data;
output egr56_valid;
input egr56_ready;
output [11:0] egr57_data;
output egr57_valid;
input egr57_ready;
output [11:0] egr58_data;
output egr58_valid;
input egr58_ready;
output [11:0] egr59_data;
output egr59_valid;
input egr59_ready;
output [11:0] egr60_data;
output egr60_valid;
input egr60_ready;
output [11:0] egr61_data;
output egr61_valid;
input egr61_ready;
output [11:0] egr62_data;
output egr62_valid;
input egr62_ready;
output [11:0] egr63_data;
output egr63_valid;
input egr63_ready;
output [11:0] egr64_data;
output egr64_valid;
input egr64_ready;
output [11:0] egr65_data;
output egr65_valid;
input egr65_ready;
output [11:0] egr66_data;
output egr66_valid;
input egr66_ready;
output [11:0] egr67_data;
output egr67_valid;
input egr67_ready;
output [11:0] egr68_data;
output egr68_valid;
input egr68_ready;
output [11:0] egr69_data;
output egr69_valid;
input egr69_ready;
output [11:0] egr70_data;
output egr70_valid;
input egr70_ready;
output [11:0] egr71_data;
output egr71_valid;
input egr71_ready;
output [11:0] egr72_data;
output egr72_valid;
input egr72_ready;
output [11:0] egr73_data;
output egr73_valid;
input egr73_ready;
output [11:0] egr74_data;
output egr74_valid;
input egr74_ready;
output [11:0] egr75_data;
output egr75_valid;
input egr75_ready;
output [11:0] egr76_data;
output egr76_valid;
input egr76_ready;
output [11:0] egr77_data;
output egr77_valid;
input egr77_ready;
output [11:0] egr78_data;
output egr78_valid;
input egr78_ready;
output [11:0] egr79_data;
output egr79_valid;
input egr79_ready;
output [11:0] egr80_data;
output egr80_valid;
input egr80_ready;
output [11:0] egr81_data;
output egr81_valid;
input egr81_ready;
output [11:0] egr82_data;
output egr82_valid;
input egr82_ready;
output [11:0] egr83_data;
output egr83_valid;
input egr83_ready;
output [11:0] egr84_data;
output egr84_valid;
input egr84_ready;
output [11:0] egr85_data;
output egr85_valid;
input egr85_ready;
output [11:0] egr86_data;
output egr86_valid;
input egr86_ready;
output [11:0] egr87_data;
output egr87_valid;
input egr87_ready;
output [11:0] egr88_data;
output egr88_valid;
input egr88_ready;
output [11:0] egr89_data;
output egr89_valid;
input egr89_ready;
output [11:0] egr90_data;
output egr90_valid;
input egr90_ready;
output [11:0] egr91_data;
output egr91_valid;
input egr91_ready;
output [11:0] egr92_data;
output egr92_valid;
input egr92_ready;
output [11:0] egr93_data;
output egr93_valid;
input egr93_ready;
output [11:0] egr94_data;
output egr94_valid;
input egr94_ready;
output [11:0] egr95_data;
output egr95_valid;
input egr95_ready;
output [11:0] egr96_data;
output egr96_valid;
input egr96_ready;
output [11:0] egr97_data;
output egr97_valid;
input egr97_ready;
output [11:0] egr98_data;
output egr98_valid;
input egr98_ready;
output [11:0] egr99_data;
output egr99_valid;
input egr99_ready;
output [11:0] egr100_data;
output egr100_valid;
input egr100_ready;
output [11:0] egr101_data;
output egr101_valid;
input egr101_ready;
output [11:0] egr102_data;
output egr102_valid;
input egr102_ready;
output [11:0] egr103_data;
output egr103_valid;
input egr103_ready;
output [11:0] egr104_data;
output egr104_valid;
input egr104_ready;
output [11:0] egr105_data;
output egr105_valid;
input egr105_ready;
output [11:0] egr106_data;
output egr106_valid;
input egr106_ready;
output [11:0] egr107_data;
output egr107_valid;
input egr107_ready;
output [11:0] egr108_data;
output egr108_valid;
input egr108_ready;
output [11:0] egr109_data;
output egr109_valid;
input egr109_ready;
output [11:0] egr110_data;
output egr110_valid;
input egr110_ready;
output [11:0] egr111_data;
output egr111_valid;
input egr111_ready;
output [11:0] egr112_data;
output egr112_valid;
input egr112_ready;
output [11:0] egr113_data;
output egr113_valid;
input egr113_ready;
output [11:0] egr114_data;
output egr114_valid;
input egr114_ready;
output [11:0] egr115_data;
output egr115_valid;
input egr115_ready;
output [11:0] egr116_data;
output egr116_valid;
input egr116_ready;
output [11:0] egr117_data;
output egr117_valid;
input egr117_ready;
output [11:0] egr118_data;
output egr118_valid;
input egr118_ready;
output [11:0] egr119_data;
output egr119_valid;
input egr119_ready;
output [11:0] egr120_data;
output egr120_valid;
input egr120_ready;
output [11:0] egr121_data;
output egr121_valid;
input egr121_ready;
output [11:0] egr122_data;
output egr122_valid;
input egr122_ready;
output [11:0] egr123_data;
output egr123_valid;
input egr123_ready;
output [11:0] egr124_data;
output egr124_valid;
input egr124_ready;
output [11:0] egr125_data;
output egr125_valid;
input egr125_ready;
output [11:0] egr126_data;
output egr126_valid;
input egr126_ready;
output [11:0] egr127_data;
output egr127_valid;
input egr127_ready;
output [11:0] egr128_data;
output egr128_valid;
input egr128_ready;
output [11:0] egr129_data;
output egr129_valid;
input egr129_ready;
output [11:0] egr130_data;
output egr130_valid;
input egr130_ready;
output [11:0] egr131_data;
output egr131_valid;
input egr131_ready;
output [11:0] egr132_data;
output egr132_valid;
input egr132_ready;
output [11:0] egr133_data;
output egr133_valid;
input egr133_ready;
output [11:0] egr134_data;
output egr134_valid;
input egr134_ready;
output [11:0] egr135_data;
output egr135_valid;
input egr135_ready;
output [11:0] egr136_data;
output egr136_valid;
input egr136_ready;
output [11:0] egr137_data;
output egr137_valid;
input egr137_ready;
output [11:0] egr138_data;
output egr138_valid;
input egr138_ready;
output [11:0] egr139_data;
output egr139_valid;
input egr139_ready;
output [11:0] egr140_data;
output egr140_valid;
input egr140_ready;
output [11:0] egr141_data;
output egr141_valid;
input egr141_ready;
output [11:0] egr142_data;
output egr142_valid;
input egr142_ready;
output [11:0] egr143_data;
output egr143_valid;
input egr143_ready;
output [11:0] egr144_data;
output egr144_valid;
input egr144_ready;
output [11:0] egr145_data;
output egr145_valid;
input egr145_ready;
output [11:0] egr146_data;
output egr146_valid;
input egr146_ready;
output [11:0] egr147_data;
output egr147_valid;
input egr147_ready;
output [11:0] egr148_data;
output egr148_valid;
input egr148_ready;
output [11:0] egr149_data;
output egr149_valid;
input egr149_ready;
output [11:0] egr150_data;
output egr150_valid;
input egr150_ready;
output [11:0] egr151_data;
output egr151_valid;
input egr151_ready;
output [11:0] egr152_data;
output egr152_valid;
input egr152_ready;
output [11:0] egr153_data;
output egr153_valid;
input egr153_ready;
output [11:0] egr154_data;
output egr154_valid;
input egr154_ready;
output [11:0] egr155_data;
output egr155_valid;
input egr155_ready;
output [11:0] egr156_data;
output egr156_valid;
input egr156_ready;
output [11:0] egr157_data;
output egr157_valid;
input egr157_ready;
output [11:0] egr158_data;
output egr158_valid;
input egr158_ready;
output [11:0] egr159_data;
output egr159_valid;
input egr159_ready;
output [11:0] egr160_data;
output egr160_valid;
input egr160_ready;
output [11:0] egr161_data;
output egr161_valid;
input egr161_ready;
output [11:0] egr162_data;
output egr162_valid;
input egr162_ready;
output [11:0] egr163_data;
output egr163_valid;
input egr163_ready;
output [11:0] egr164_data;
output egr164_valid;
input egr164_ready;
output [11:0] egr165_data;
output egr165_valid;
input egr165_ready;
output [11:0] egr166_data;
output egr166_valid;
input egr166_ready;
output [11:0] egr167_data;
output egr167_valid;
input egr167_ready;
output [11:0] egr168_data;
output egr168_valid;
input egr168_ready;
output [11:0] egr169_data;
output egr169_valid;
input egr169_ready;
output [11:0] egr170_data;
output egr170_valid;
input egr170_ready;
output [11:0] egr171_data;
output egr171_valid;
input egr171_ready;
output [11:0] egr172_data;
output egr172_valid;
input egr172_ready;
output [11:0] egr173_data;
output egr173_valid;
input egr173_ready;
output [11:0] egr174_data;
output egr174_valid;
input egr174_ready;
output [11:0] egr175_data;
output egr175_valid;
input egr175_ready;
output [11:0] egr176_data;
output egr176_valid;
input egr176_ready;
output [11:0] egr177_data;
output egr177_valid;
input egr177_ready;
output [11:0] egr178_data;
output egr178_valid;
input egr178_ready;
output [11:0] egr179_data;
output egr179_valid;
input egr179_ready;
output [11:0] egr180_data;
output egr180_valid;
input egr180_ready;
output [11:0] egr181_data;
output egr181_valid;
input egr181_ready;
output [11:0] egr182_data;
output egr182_valid;
input egr182_ready;
output [11:0] egr183_data;
output egr183_valid;
input egr183_ready;
output [11:0] egr184_data;
output egr184_valid;
input egr184_ready;
output [11:0] egr185_data;
output egr185_valid;
input egr185_ready;
output [11:0] egr186_data;
output egr186_valid;
input egr186_ready;
output [11:0] egr187_data;
output egr187_valid;
input egr187_ready;
output [11:0] egr188_data;
output egr188_valid;
input egr188_ready;
output [11:0] egr189_data;
output egr189_valid;
input egr189_ready;
output [11:0] egr190_data;
output egr190_valid;
input egr190_ready;
output [11:0] egr191_data;
output egr191_valid;
input egr191_ready;
output [11:0] egr192_data;
output egr192_valid;
input egr192_ready;
output [11:0] egr193_data;
output egr193_valid;
input egr193_ready;
output [11:0] egr194_data;
output egr194_valid;
input egr194_ready;
output [11:0] egr195_data;
output egr195_valid;
input egr195_ready;
output [11:0] egr196_data;
output egr196_valid;
input egr196_ready;
output [11:0] egr197_data;
output egr197_valid;
input egr197_ready;
output [11:0] egr198_data;
output egr198_valid;
input egr198_ready;
output [11:0] egr199_data;
output egr199_valid;
input egr199_ready;
output [11:0] egr200_data;
output egr200_valid;
input egr200_ready;
output [11:0] egr201_data;
output egr201_valid;
input egr201_ready;
output [11:0] egr202_data;
output egr202_valid;
input egr202_ready;
output [11:0] egr203_data;
output egr203_valid;
input egr203_ready;
output [11:0] egr204_data;
output egr204_valid;
input egr204_ready;
output [11:0] egr205_data;
output egr205_valid;
input egr205_ready;
output [11:0] egr206_data;
output egr206_valid;
input egr206_ready;
output [11:0] egr207_data;
output egr207_valid;
input egr207_ready;
output [11:0] egr208_data;
output egr208_valid;
input egr208_ready;
output [11:0] egr209_data;
output egr209_valid;
input egr209_ready;
output [11:0] egr210_data;
output egr210_valid;
input egr210_ready;
output [11:0] egr211_data;
output egr211_valid;
input egr211_ready;
output [11:0] egr212_data;
output egr212_valid;
input egr212_ready;
output [11:0] egr213_data;
output egr213_valid;
input egr213_ready;
output [11:0] egr214_data;
output egr214_valid;
input egr214_ready;
output [11:0] egr215_data;
output egr215_valid;
input egr215_ready;
output [11:0] egr216_data;
output egr216_valid;
input egr216_ready;
output [11:0] egr217_data;
output egr217_valid;
input egr217_ready;
output [11:0] egr218_data;
output egr218_valid;
input egr218_ready;
output [11:0] egr219_data;
output egr219_valid;
input egr219_ready;
output [11:0] egr220_data;
output egr220_valid;
input egr220_ready;
output [11:0] egr221_data;
output egr221_valid;
input egr221_ready;
output [11:0] egr222_data;
output egr222_valid;
input egr222_ready;
output [11:0] egr223_data;
output egr223_valid;
input egr223_ready;
output [11:0] egr224_data;
output egr224_valid;
input egr224_ready;
output [11:0] egr225_data;
output egr225_valid;
input egr225_ready;
output [11:0] egr226_data;
output egr226_valid;
input egr226_ready;
output [11:0] egr227_data;
output egr227_valid;
input egr227_ready;
output [11:0] egr228_data;
output egr228_valid;
input egr228_ready;
output [11:0] egr229_data;
output egr229_valid;
input egr229_ready;
output [11:0] egr230_data;
output egr230_valid;
input egr230_ready;
output [11:0] egr231_data;
output egr231_valid;
input egr231_ready;
output [11:0] egr232_data;
output egr232_valid;
input egr232_ready;
output [11:0] egr233_data;
output egr233_valid;
input egr233_ready;
output [11:0] egr234_data;
output egr234_valid;
input egr234_ready;
output [11:0] egr235_data;
output egr235_valid;
input egr235_ready;
output [11:0] egr236_data;
output egr236_valid;
input egr236_ready;
output [11:0] egr237_data;
output egr237_valid;
input egr237_ready;
output [11:0] egr238_data;
output egr238_valid;
input egr238_ready;
output [11:0] egr239_data;
output egr239_valid;
input egr239_ready;
output [11:0] egr240_data;
output egr240_valid;
input egr240_ready;
output [11:0] egr241_data;
output egr241_valid;
input egr241_ready;
output [11:0] egr242_data;
output egr242_valid;
input egr242_ready;
output [11:0] egr243_data;
output egr243_valid;
input egr243_ready;
output [11:0] egr244_data;
output egr244_valid;
input egr244_ready;
output [11:0] egr245_data;
output egr245_valid;
input egr245_ready;
output [11:0] egr246_data;
output egr246_valid;
input egr246_ready;
output [11:0] egr247_data;
output egr247_valid;
input egr247_ready;
output [11:0] egr248_data;
output egr248_valid;
input egr248_ready;
output [11:0] egr249_data;
output egr249_valid;
input egr249_ready;
output [11:0] egr250_data;
output egr250_valid;
input egr250_ready;
output [11:0] egr251_data;
output egr251_valid;
input egr251_ready;
output [11:0] egr252_data;
output egr252_valid;
input egr252_ready;
output [11:0] egr253_data;
output egr253_valid;
input egr253_ready;
output [11:0] egr254_data;
output egr254_valid;
input egr254_ready;
output [11:0] egr255_data;
output egr255_valid;
input egr255_ready;
output [11:0] egr256_data;
output egr256_valid;
input egr256_ready;
output [11:0] egr257_data;
output egr257_valid;
input egr257_ready;


// Ingress and Egress are short circuited based on condition


wire assign egress0_ds_pkt       = (demux_select== 9'd0) ? ingress_ds_pkt       : 9'd0;
wire assign egress1_ds_pkt       = (demux_select== 9'd1) ? ingress_ds_pkt       : 9'd0;
wire assign egress2_ds_pkt       = (demux_select== 9'd2) ? ingress_ds_pkt       : 9'd0;
wire assign egress3_ds_pkt       = (demux_select== 9'd3) ? ingress_ds_pkt       : 9'd0;
wire assign egress4_ds_pkt       = (demux_select== 9'd4) ? ingress_ds_pkt       : 9'd0;
wire assign egress5_ds_pkt       = (demux_select== 9'd5) ? ingress_ds_pkt       : 9'd0;
wire assign egress6_ds_pkt       = (demux_select== 9'd6) ? ingress_ds_pkt       : 9'd0;
wire assign egress7_ds_pkt       = (demux_select== 9'd7) ? ingress_ds_pkt       : 9'd0;
wire assign egress8_ds_pkt       = (demux_select== 9'd8) ? ingress_ds_pkt       : 9'd0;
wire assign egress9_ds_pkt       = (demux_select== 9'd9) ? ingress_ds_pkt       : 9'd0;
wire assign egress10_ds_pkt       = (demux_select== 9'd10) ? ingress_ds_pkt       : 9'd0;
wire assign egress11_ds_pkt       = (demux_select== 9'd11) ? ingress_ds_pkt       : 9'd0;
wire assign egress12_ds_pkt       = (demux_select== 9'd12) ? ingress_ds_pkt       : 9'd0;
wire assign egress13_ds_pkt       = (demux_select== 9'd13) ? ingress_ds_pkt       : 9'd0;
wire assign egress14_ds_pkt       = (demux_select== 9'd14) ? ingress_ds_pkt       : 9'd0;
wire assign egress15_ds_pkt       = (demux_select== 9'd15) ? ingress_ds_pkt       : 9'd0;
wire assign egress16_ds_pkt       = (demux_select== 9'd16) ? ingress_ds_pkt       : 9'd0;
wire assign egress17_ds_pkt       = (demux_select== 9'd17) ? ingress_ds_pkt       : 9'd0;
wire assign egress18_ds_pkt       = (demux_select== 9'd18) ? ingress_ds_pkt       : 9'd0;
wire assign egress19_ds_pkt       = (demux_select== 9'd19) ? ingress_ds_pkt       : 9'd0;
wire assign egress20_ds_pkt       = (demux_select== 9'd20) ? ingress_ds_pkt       : 9'd0;
wire assign egress21_ds_pkt       = (demux_select== 9'd21) ? ingress_ds_pkt       : 9'd0;
wire assign egress22_ds_pkt       = (demux_select== 9'd22) ? ingress_ds_pkt       : 9'd0;
wire assign egress23_ds_pkt       = (demux_select== 9'd23) ? ingress_ds_pkt       : 9'd0;
wire assign egress24_ds_pkt       = (demux_select== 9'd24) ? ingress_ds_pkt       : 9'd0;
wire assign egress25_ds_pkt       = (demux_select== 9'd25) ? ingress_ds_pkt       : 9'd0;
wire assign egress26_ds_pkt       = (demux_select== 9'd26) ? ingress_ds_pkt       : 9'd0;
wire assign egress27_ds_pkt       = (demux_select== 9'd27) ? ingress_ds_pkt       : 9'd0;
wire assign egress28_ds_pkt       = (demux_select== 9'd28) ? ingress_ds_pkt       : 9'd0;
wire assign egress29_ds_pkt       = (demux_select== 9'd29) ? ingress_ds_pkt       : 9'd0;
wire assign egress30_ds_pkt       = (demux_select== 9'd30) ? ingress_ds_pkt       : 9'd0;
wire assign egress31_ds_pkt       = (demux_select== 9'd31) ? ingress_ds_pkt       : 9'd0;
wire assign egress32_ds_pkt       = (demux_select== 9'd32) ? ingress_ds_pkt       : 9'd0;
wire assign egress33_ds_pkt       = (demux_select== 9'd33) ? ingress_ds_pkt       : 9'd0;
wire assign egress34_ds_pkt       = (demux_select== 9'd34) ? ingress_ds_pkt       : 9'd0;
wire assign egress35_ds_pkt       = (demux_select== 9'd35) ? ingress_ds_pkt       : 9'd0;
wire assign egress36_ds_pkt       = (demux_select== 9'd36) ? ingress_ds_pkt       : 9'd0;
wire assign egress37_ds_pkt       = (demux_select== 9'd37) ? ingress_ds_pkt       : 9'd0;
wire assign egress38_ds_pkt       = (demux_select== 9'd38) ? ingress_ds_pkt       : 9'd0;
wire assign egress39_ds_pkt       = (demux_select== 9'd39) ? ingress_ds_pkt       : 9'd0;
wire assign egress40_ds_pkt       = (demux_select== 9'd40) ? ingress_ds_pkt       : 9'd0;
wire assign egress41_ds_pkt       = (demux_select== 9'd41) ? ingress_ds_pkt       : 9'd0;
wire assign egress42_ds_pkt       = (demux_select== 9'd42) ? ingress_ds_pkt       : 9'd0;
wire assign egress43_ds_pkt       = (demux_select== 9'd43) ? ingress_ds_pkt       : 9'd0;
wire assign egress44_ds_pkt       = (demux_select== 9'd44) ? ingress_ds_pkt       : 9'd0;
wire assign egress45_ds_pkt       = (demux_select== 9'd45) ? ingress_ds_pkt       : 9'd0;
wire assign egress46_ds_pkt       = (demux_select== 9'd46) ? ingress_ds_pkt       : 9'd0;
wire assign egress47_ds_pkt       = (demux_select== 9'd47) ? ingress_ds_pkt       : 9'd0;
wire assign egress48_ds_pkt       = (demux_select== 9'd48) ? ingress_ds_pkt       : 9'd0;
wire assign egress49_ds_pkt       = (demux_select== 9'd49) ? ingress_ds_pkt       : 9'd0;
wire assign egress50_ds_pkt       = (demux_select== 9'd50) ? ingress_ds_pkt       : 9'd0;
wire assign egress51_ds_pkt       = (demux_select== 9'd51) ? ingress_ds_pkt       : 9'd0;
wire assign egress52_ds_pkt       = (demux_select== 9'd52) ? ingress_ds_pkt       : 9'd0;
wire assign egress53_ds_pkt       = (demux_select== 9'd53) ? ingress_ds_pkt       : 9'd0;
wire assign egress54_ds_pkt       = (demux_select== 9'd54) ? ingress_ds_pkt       : 9'd0;
wire assign egress55_ds_pkt       = (demux_select== 9'd55) ? ingress_ds_pkt       : 9'd0;
wire assign egress56_ds_pkt       = (demux_select== 9'd56) ? ingress_ds_pkt       : 9'd0;
wire assign egress57_ds_pkt       = (demux_select== 9'd57) ? ingress_ds_pkt       : 9'd0;
wire assign egress58_ds_pkt       = (demux_select== 9'd58) ? ingress_ds_pkt       : 9'd0;
wire assign egress59_ds_pkt       = (demux_select== 9'd59) ? ingress_ds_pkt       : 9'd0;
wire assign egress60_ds_pkt       = (demux_select== 9'd60) ? ingress_ds_pkt       : 9'd0;
wire assign egress61_ds_pkt       = (demux_select== 9'd61) ? ingress_ds_pkt       : 9'd0;
wire assign egress62_ds_pkt       = (demux_select== 9'd62) ? ingress_ds_pkt       : 9'd0;
wire assign egress63_ds_pkt       = (demux_select== 9'd63) ? ingress_ds_pkt       : 9'd0;
wire assign egress64_ds_pkt       = (demux_select== 9'd64) ? ingress_ds_pkt       : 9'd0;
wire assign egress65_ds_pkt       = (demux_select== 9'd65) ? ingress_ds_pkt       : 9'd0;
wire assign egress66_ds_pkt       = (demux_select== 9'd66) ? ingress_ds_pkt       : 9'd0;
wire assign egress67_ds_pkt       = (demux_select== 9'd67) ? ingress_ds_pkt       : 9'd0;
wire assign egress68_ds_pkt       = (demux_select== 9'd68) ? ingress_ds_pkt       : 9'd0;
wire assign egress69_ds_pkt       = (demux_select== 9'd69) ? ingress_ds_pkt       : 9'd0;
wire assign egress70_ds_pkt       = (demux_select== 9'd70) ? ingress_ds_pkt       : 9'd0;
wire assign egress71_ds_pkt       = (demux_select== 9'd71) ? ingress_ds_pkt       : 9'd0;
wire assign egress72_ds_pkt       = (demux_select== 9'd72) ? ingress_ds_pkt       : 9'd0;
wire assign egress73_ds_pkt       = (demux_select== 9'd73) ? ingress_ds_pkt       : 9'd0;
wire assign egress74_ds_pkt       = (demux_select== 9'd74) ? ingress_ds_pkt       : 9'd0;
wire assign egress75_ds_pkt       = (demux_select== 9'd75) ? ingress_ds_pkt       : 9'd0;
wire assign egress76_ds_pkt       = (demux_select== 9'd76) ? ingress_ds_pkt       : 9'd0;
wire assign egress77_ds_pkt       = (demux_select== 9'd77) ? ingress_ds_pkt       : 9'd0;
wire assign egress78_ds_pkt       = (demux_select== 9'd78) ? ingress_ds_pkt       : 9'd0;
wire assign egress79_ds_pkt       = (demux_select== 9'd79) ? ingress_ds_pkt       : 9'd0;
wire assign egress80_ds_pkt       = (demux_select== 9'd80) ? ingress_ds_pkt       : 9'd0;
wire assign egress81_ds_pkt       = (demux_select== 9'd81) ? ingress_ds_pkt       : 9'd0;
wire assign egress82_ds_pkt       = (demux_select== 9'd82) ? ingress_ds_pkt       : 9'd0;
wire assign egress83_ds_pkt       = (demux_select== 9'd83) ? ingress_ds_pkt       : 9'd0;
wire assign egress84_ds_pkt       = (demux_select== 9'd84) ? ingress_ds_pkt       : 9'd0;
wire assign egress85_ds_pkt       = (demux_select== 9'd85) ? ingress_ds_pkt       : 9'd0;
wire assign egress86_ds_pkt       = (demux_select== 9'd86) ? ingress_ds_pkt       : 9'd0;
wire assign egress87_ds_pkt       = (demux_select== 9'd87) ? ingress_ds_pkt       : 9'd0;
wire assign egress88_ds_pkt       = (demux_select== 9'd88) ? ingress_ds_pkt       : 9'd0;
wire assign egress89_ds_pkt       = (demux_select== 9'd89) ? ingress_ds_pkt       : 9'd0;
wire assign egress90_ds_pkt       = (demux_select== 9'd90) ? ingress_ds_pkt       : 9'd0;
wire assign egress91_ds_pkt       = (demux_select== 9'd91) ? ingress_ds_pkt       : 9'd0;
wire assign egress92_ds_pkt       = (demux_select== 9'd92) ? ingress_ds_pkt       : 9'd0;
wire assign egress93_ds_pkt       = (demux_select== 9'd93) ? ingress_ds_pkt       : 9'd0;
wire assign egress94_ds_pkt       = (demux_select== 9'd94) ? ingress_ds_pkt       : 9'd0;
wire assign egress95_ds_pkt       = (demux_select== 9'd95) ? ingress_ds_pkt       : 9'd0;
wire assign egress96_ds_pkt       = (demux_select== 9'd96) ? ingress_ds_pkt       : 9'd0;
wire assign egress97_ds_pkt       = (demux_select== 9'd97) ? ingress_ds_pkt       : 9'd0;
wire assign egress98_ds_pkt       = (demux_select== 9'd98) ? ingress_ds_pkt       : 9'd0;
wire assign egress99_ds_pkt       = (demux_select== 9'd99) ? ingress_ds_pkt       : 9'd0;
wire assign egress100_ds_pkt       = (demux_select== 9'd100) ? ingress_ds_pkt       : 9'd0;
wire assign egress101_ds_pkt       = (demux_select== 9'd101) ? ingress_ds_pkt       : 9'd0;
wire assign egress102_ds_pkt       = (demux_select== 9'd102) ? ingress_ds_pkt       : 9'd0;
wire assign egress103_ds_pkt       = (demux_select== 9'd103) ? ingress_ds_pkt       : 9'd0;
wire assign egress104_ds_pkt       = (demux_select== 9'd104) ? ingress_ds_pkt       : 9'd0;
wire assign egress105_ds_pkt       = (demux_select== 9'd105) ? ingress_ds_pkt       : 9'd0;
wire assign egress106_ds_pkt       = (demux_select== 9'd106) ? ingress_ds_pkt       : 9'd0;
wire assign egress107_ds_pkt       = (demux_select== 9'd107) ? ingress_ds_pkt       : 9'd0;
wire assign egress108_ds_pkt       = (demux_select== 9'd108) ? ingress_ds_pkt       : 9'd0;
wire assign egress109_ds_pkt       = (demux_select== 9'd109) ? ingress_ds_pkt       : 9'd0;
wire assign egress110_ds_pkt       = (demux_select== 9'd110) ? ingress_ds_pkt       : 9'd0;
wire assign egress111_ds_pkt       = (demux_select== 9'd111) ? ingress_ds_pkt       : 9'd0;
wire assign egress112_ds_pkt       = (demux_select== 9'd112) ? ingress_ds_pkt       : 9'd0;
wire assign egress113_ds_pkt       = (demux_select== 9'd113) ? ingress_ds_pkt       : 9'd0;
wire assign egress114_ds_pkt       = (demux_select== 9'd114) ? ingress_ds_pkt       : 9'd0;
wire assign egress115_ds_pkt       = (demux_select== 9'd115) ? ingress_ds_pkt       : 9'd0;
wire assign egress116_ds_pkt       = (demux_select== 9'd116) ? ingress_ds_pkt       : 9'd0;
wire assign egress117_ds_pkt       = (demux_select== 9'd117) ? ingress_ds_pkt       : 9'd0;
wire assign egress118_ds_pkt       = (demux_select== 9'd118) ? ingress_ds_pkt       : 9'd0;
wire assign egress119_ds_pkt       = (demux_select== 9'd119) ? ingress_ds_pkt       : 9'd0;
wire assign egress120_ds_pkt       = (demux_select== 9'd120) ? ingress_ds_pkt       : 9'd0;
wire assign egress121_ds_pkt       = (demux_select== 9'd121) ? ingress_ds_pkt       : 9'd0;
wire assign egress122_ds_pkt       = (demux_select== 9'd122) ? ingress_ds_pkt       : 9'd0;
wire assign egress123_ds_pkt       = (demux_select== 9'd123) ? ingress_ds_pkt       : 9'd0;
wire assign egress124_ds_pkt       = (demux_select== 9'd124) ? ingress_ds_pkt       : 9'd0;
wire assign egress125_ds_pkt       = (demux_select== 9'd125) ? ingress_ds_pkt       : 9'd0;
wire assign egress126_ds_pkt       = (demux_select== 9'd126) ? ingress_ds_pkt       : 9'd0;
wire assign egress127_ds_pkt       = (demux_select== 9'd127) ? ingress_ds_pkt       : 9'd0;
wire assign egress128_ds_pkt       = (demux_select== 9'd128) ? ingress_ds_pkt       : 9'd0;
wire assign egress129_ds_pkt       = (demux_select== 9'd129) ? ingress_ds_pkt       : 9'd0;
wire assign egress130_ds_pkt       = (demux_select== 9'd130) ? ingress_ds_pkt       : 9'd0;
wire assign egress131_ds_pkt       = (demux_select== 9'd131) ? ingress_ds_pkt       : 9'd0;
wire assign egress132_ds_pkt       = (demux_select== 9'd132) ? ingress_ds_pkt       : 9'd0;
wire assign egress133_ds_pkt       = (demux_select== 9'd133) ? ingress_ds_pkt       : 9'd0;
wire assign egress134_ds_pkt       = (demux_select== 9'd134) ? ingress_ds_pkt       : 9'd0;
wire assign egress135_ds_pkt       = (demux_select== 9'd135) ? ingress_ds_pkt       : 9'd0;
wire assign egress136_ds_pkt       = (demux_select== 9'd136) ? ingress_ds_pkt       : 9'd0;
wire assign egress137_ds_pkt       = (demux_select== 9'd137) ? ingress_ds_pkt       : 9'd0;
wire assign egress138_ds_pkt       = (demux_select== 9'd138) ? ingress_ds_pkt       : 9'd0;
wire assign egress139_ds_pkt       = (demux_select== 9'd139) ? ingress_ds_pkt       : 9'd0;
wire assign egress140_ds_pkt       = (demux_select== 9'd140) ? ingress_ds_pkt       : 9'd0;
wire assign egress141_ds_pkt       = (demux_select== 9'd141) ? ingress_ds_pkt       : 9'd0;
wire assign egress142_ds_pkt       = (demux_select== 9'd142) ? ingress_ds_pkt       : 9'd0;
wire assign egress143_ds_pkt       = (demux_select== 9'd143) ? ingress_ds_pkt       : 9'd0;
wire assign egress144_ds_pkt       = (demux_select== 9'd144) ? ingress_ds_pkt       : 9'd0;
wire assign egress145_ds_pkt       = (demux_select== 9'd145) ? ingress_ds_pkt       : 9'd0;
wire assign egress146_ds_pkt       = (demux_select== 9'd146) ? ingress_ds_pkt       : 9'd0;
wire assign egress147_ds_pkt       = (demux_select== 9'd147) ? ingress_ds_pkt       : 9'd0;
wire assign egress148_ds_pkt       = (demux_select== 9'd148) ? ingress_ds_pkt       : 9'd0;
wire assign egress149_ds_pkt       = (demux_select== 9'd149) ? ingress_ds_pkt       : 9'd0;
wire assign egress150_ds_pkt       = (demux_select== 9'd150) ? ingress_ds_pkt       : 9'd0;
wire assign egress151_ds_pkt       = (demux_select== 9'd151) ? ingress_ds_pkt       : 9'd0;
wire assign egress152_ds_pkt       = (demux_select== 9'd152) ? ingress_ds_pkt       : 9'd0;
wire assign egress153_ds_pkt       = (demux_select== 9'd153) ? ingress_ds_pkt       : 9'd0;
wire assign egress154_ds_pkt       = (demux_select== 9'd154) ? ingress_ds_pkt       : 9'd0;
wire assign egress155_ds_pkt       = (demux_select== 9'd155) ? ingress_ds_pkt       : 9'd0;
wire assign egress156_ds_pkt       = (demux_select== 9'd156) ? ingress_ds_pkt       : 9'd0;
wire assign egress157_ds_pkt       = (demux_select== 9'd157) ? ingress_ds_pkt       : 9'd0;
wire assign egress158_ds_pkt       = (demux_select== 9'd158) ? ingress_ds_pkt       : 9'd0;
wire assign egress159_ds_pkt       = (demux_select== 9'd159) ? ingress_ds_pkt       : 9'd0;
wire assign egress160_ds_pkt       = (demux_select== 9'd160) ? ingress_ds_pkt       : 9'd0;
wire assign egress161_ds_pkt       = (demux_select== 9'd161) ? ingress_ds_pkt       : 9'd0;
wire assign egress162_ds_pkt       = (demux_select== 9'd162) ? ingress_ds_pkt       : 9'd0;
wire assign egress163_ds_pkt       = (demux_select== 9'd163) ? ingress_ds_pkt       : 9'd0;
wire assign egress164_ds_pkt       = (demux_select== 9'd164) ? ingress_ds_pkt       : 9'd0;
wire assign egress165_ds_pkt       = (demux_select== 9'd165) ? ingress_ds_pkt       : 9'd0;
wire assign egress166_ds_pkt       = (demux_select== 9'd166) ? ingress_ds_pkt       : 9'd0;
wire assign egress167_ds_pkt       = (demux_select== 9'd167) ? ingress_ds_pkt       : 9'd0;
wire assign egress168_ds_pkt       = (demux_select== 9'd168) ? ingress_ds_pkt       : 9'd0;
wire assign egress169_ds_pkt       = (demux_select== 9'd169) ? ingress_ds_pkt       : 9'd0;
wire assign egress170_ds_pkt       = (demux_select== 9'd170) ? ingress_ds_pkt       : 9'd0;
wire assign egress171_ds_pkt       = (demux_select== 9'd171) ? ingress_ds_pkt       : 9'd0;
wire assign egress172_ds_pkt       = (demux_select== 9'd172) ? ingress_ds_pkt       : 9'd0;
wire assign egress173_ds_pkt       = (demux_select== 9'd173) ? ingress_ds_pkt       : 9'd0;
wire assign egress174_ds_pkt       = (demux_select== 9'd174) ? ingress_ds_pkt       : 9'd0;
wire assign egress175_ds_pkt       = (demux_select== 9'd175) ? ingress_ds_pkt       : 9'd0;
wire assign egress176_ds_pkt       = (demux_select== 9'd176) ? ingress_ds_pkt       : 9'd0;
wire assign egress177_ds_pkt       = (demux_select== 9'd177) ? ingress_ds_pkt       : 9'd0;
wire assign egress178_ds_pkt       = (demux_select== 9'd178) ? ingress_ds_pkt       : 9'd0;
wire assign egress179_ds_pkt       = (demux_select== 9'd179) ? ingress_ds_pkt       : 9'd0;
wire assign egress180_ds_pkt       = (demux_select== 9'd180) ? ingress_ds_pkt       : 9'd0;
wire assign egress181_ds_pkt       = (demux_select== 9'd181) ? ingress_ds_pkt       : 9'd0;
wire assign egress182_ds_pkt       = (demux_select== 9'd182) ? ingress_ds_pkt       : 9'd0;
wire assign egress183_ds_pkt       = (demux_select== 9'd183) ? ingress_ds_pkt       : 9'd0;
wire assign egress184_ds_pkt       = (demux_select== 9'd184) ? ingress_ds_pkt       : 9'd0;
wire assign egress185_ds_pkt       = (demux_select== 9'd185) ? ingress_ds_pkt       : 9'd0;
wire assign egress186_ds_pkt       = (demux_select== 9'd186) ? ingress_ds_pkt       : 9'd0;
wire assign egress187_ds_pkt       = (demux_select== 9'd187) ? ingress_ds_pkt       : 9'd0;
wire assign egress188_ds_pkt       = (demux_select== 9'd188) ? ingress_ds_pkt       : 9'd0;
wire assign egress189_ds_pkt       = (demux_select== 9'd189) ? ingress_ds_pkt       : 9'd0;
wire assign egress190_ds_pkt       = (demux_select== 9'd190) ? ingress_ds_pkt       : 9'd0;
wire assign egress191_ds_pkt       = (demux_select== 9'd191) ? ingress_ds_pkt       : 9'd0;
wire assign egress192_ds_pkt       = (demux_select== 9'd192) ? ingress_ds_pkt       : 9'd0;
wire assign egress193_ds_pkt       = (demux_select== 9'd193) ? ingress_ds_pkt       : 9'd0;
wire assign egress194_ds_pkt       = (demux_select== 9'd194) ? ingress_ds_pkt       : 9'd0;
wire assign egress195_ds_pkt       = (demux_select== 9'd195) ? ingress_ds_pkt       : 9'd0;
wire assign egress196_ds_pkt       = (demux_select== 9'd196) ? ingress_ds_pkt       : 9'd0;
wire assign egress197_ds_pkt       = (demux_select== 9'd197) ? ingress_ds_pkt       : 9'd0;
wire assign egress198_ds_pkt       = (demux_select== 9'd198) ? ingress_ds_pkt       : 9'd0;
wire assign egress199_ds_pkt       = (demux_select== 9'd199) ? ingress_ds_pkt       : 9'd0;
wire assign egress200_ds_pkt       = (demux_select== 9'd200) ? ingress_ds_pkt       : 9'd0;
wire assign egress201_ds_pkt       = (demux_select== 9'd201) ? ingress_ds_pkt       : 9'd0;
wire assign egress202_ds_pkt       = (demux_select== 9'd202) ? ingress_ds_pkt       : 9'd0;
wire assign egress203_ds_pkt       = (demux_select== 9'd203) ? ingress_ds_pkt       : 9'd0;
wire assign egress204_ds_pkt       = (demux_select== 9'd204) ? ingress_ds_pkt       : 9'd0;
wire assign egress205_ds_pkt       = (demux_select== 9'd205) ? ingress_ds_pkt       : 9'd0;
wire assign egress206_ds_pkt       = (demux_select== 9'd206) ? ingress_ds_pkt       : 9'd0;
wire assign egress207_ds_pkt       = (demux_select== 9'd207) ? ingress_ds_pkt       : 9'd0;
wire assign egress208_ds_pkt       = (demux_select== 9'd208) ? ingress_ds_pkt       : 9'd0;
wire assign egress209_ds_pkt       = (demux_select== 9'd209) ? ingress_ds_pkt       : 9'd0;
wire assign egress210_ds_pkt       = (demux_select== 9'd210) ? ingress_ds_pkt       : 9'd0;
wire assign egress211_ds_pkt       = (demux_select== 9'd211) ? ingress_ds_pkt       : 9'd0;
wire assign egress212_ds_pkt       = (demux_select== 9'd212) ? ingress_ds_pkt       : 9'd0;
wire assign egress213_ds_pkt       = (demux_select== 9'd213) ? ingress_ds_pkt       : 9'd0;
wire assign egress214_ds_pkt       = (demux_select== 9'd214) ? ingress_ds_pkt       : 9'd0;
wire assign egress215_ds_pkt       = (demux_select== 9'd215) ? ingress_ds_pkt       : 9'd0;
wire assign egress216_ds_pkt       = (demux_select== 9'd216) ? ingress_ds_pkt       : 9'd0;
wire assign egress217_ds_pkt       = (demux_select== 9'd217) ? ingress_ds_pkt       : 9'd0;
wire assign egress218_ds_pkt       = (demux_select== 9'd218) ? ingress_ds_pkt       : 9'd0;
wire assign egress219_ds_pkt       = (demux_select== 9'd219) ? ingress_ds_pkt       : 9'd0;
wire assign egress220_ds_pkt       = (demux_select== 9'd220) ? ingress_ds_pkt       : 9'd0;
wire assign egress221_ds_pkt       = (demux_select== 9'd221) ? ingress_ds_pkt       : 9'd0;
wire assign egress222_ds_pkt       = (demux_select== 9'd222) ? ingress_ds_pkt       : 9'd0;
wire assign egress223_ds_pkt       = (demux_select== 9'd223) ? ingress_ds_pkt       : 9'd0;
wire assign egress224_ds_pkt       = (demux_select== 9'd224) ? ingress_ds_pkt       : 9'd0;
wire assign egress225_ds_pkt       = (demux_select== 9'd225) ? ingress_ds_pkt       : 9'd0;
wire assign egress226_ds_pkt       = (demux_select== 9'd226) ? ingress_ds_pkt       : 9'd0;
wire assign egress227_ds_pkt       = (demux_select== 9'd227) ? ingress_ds_pkt       : 9'd0;
wire assign egress228_ds_pkt       = (demux_select== 9'd228) ? ingress_ds_pkt       : 9'd0;
wire assign egress229_ds_pkt       = (demux_select== 9'd229) ? ingress_ds_pkt       : 9'd0;
wire assign egress230_ds_pkt       = (demux_select== 9'd230) ? ingress_ds_pkt       : 9'd0;
wire assign egress231_ds_pkt       = (demux_select== 9'd231) ? ingress_ds_pkt       : 9'd0;
wire assign egress232_ds_pkt       = (demux_select== 9'd232) ? ingress_ds_pkt       : 9'd0;
wire assign egress233_ds_pkt       = (demux_select== 9'd233) ? ingress_ds_pkt       : 9'd0;
wire assign egress234_ds_pkt       = (demux_select== 9'd234) ? ingress_ds_pkt       : 9'd0;
wire assign egress235_ds_pkt       = (demux_select== 9'd235) ? ingress_ds_pkt       : 9'd0;
wire assign egress236_ds_pkt       = (demux_select== 9'd236) ? ingress_ds_pkt       : 9'd0;
wire assign egress237_ds_pkt       = (demux_select== 9'd237) ? ingress_ds_pkt       : 9'd0;
wire assign egress238_ds_pkt       = (demux_select== 9'd238) ? ingress_ds_pkt       : 9'd0;
wire assign egress239_ds_pkt       = (demux_select== 9'd239) ? ingress_ds_pkt       : 9'd0;
wire assign egress240_ds_pkt       = (demux_select== 9'd240) ? ingress_ds_pkt       : 9'd0;
wire assign egress241_ds_pkt       = (demux_select== 9'd241) ? ingress_ds_pkt       : 9'd0;
wire assign egress242_ds_pkt       = (demux_select== 9'd242) ? ingress_ds_pkt       : 9'd0;
wire assign egress243_ds_pkt       = (demux_select== 9'd243) ? ingress_ds_pkt       : 9'd0;
wire assign egress244_ds_pkt       = (demux_select== 9'd244) ? ingress_ds_pkt       : 9'd0;
wire assign egress245_ds_pkt       = (demux_select== 9'd245) ? ingress_ds_pkt       : 9'd0;
wire assign egress246_ds_pkt       = (demux_select== 9'd246) ? ingress_ds_pkt       : 9'd0;
wire assign egress247_ds_pkt       = (demux_select== 9'd247) ? ingress_ds_pkt       : 9'd0;
wire assign egress248_ds_pkt       = (demux_select== 9'd248) ? ingress_ds_pkt       : 9'd0;
wire assign egress249_ds_pkt       = (demux_select== 9'd249) ? ingress_ds_pkt       : 9'd0;
wire assign egress250_ds_pkt       = (demux_select== 9'd250) ? ingress_ds_pkt       : 9'd0;
wire assign egress251_ds_pkt       = (demux_select== 9'd251) ? ingress_ds_pkt       : 9'd0;
wire assign egress252_ds_pkt       = (demux_select== 9'd252) ? ingress_ds_pkt       : 9'd0;
wire assign egress253_ds_pkt       = (demux_select== 9'd253) ? ingress_ds_pkt       : 9'd0;
wire assign egress254_ds_pkt       = (demux_select== 9'd254) ? ingress_ds_pkt       : 9'd0;
wire assign egress255_ds_pkt       = (demux_select== 9'd255) ? ingress_ds_pkt       : 9'd0;
wire assign egress256_ds_pkt       = (demux_select== 9'd256) ? ingress_ds_pkt       : 9'd0;
wire assign egress257_ds_pkt       = (demux_select== 9'd257) ? ingress_ds_pkt       : 9'd0;
wire assign egress0_ds_pkt_valid = (demux_select== 9'd0) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress1_ds_pkt_valid = (demux_select== 9'd1) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress2_ds_pkt_valid = (demux_select== 9'd2) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress3_ds_pkt_valid = (demux_select== 9'd3) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress4_ds_pkt_valid = (demux_select== 9'd4) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress5_ds_pkt_valid = (demux_select== 9'd5) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress6_ds_pkt_valid = (demux_select== 9'd6) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress7_ds_pkt_valid = (demux_select== 9'd7) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress8_ds_pkt_valid = (demux_select== 9'd8) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress9_ds_pkt_valid = (demux_select== 9'd9) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress10_ds_pkt_valid = (demux_select== 9'd10) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress11_ds_pkt_valid = (demux_select== 9'd11) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress12_ds_pkt_valid = (demux_select== 9'd12) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress13_ds_pkt_valid = (demux_select== 9'd13) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress14_ds_pkt_valid = (demux_select== 9'd14) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress15_ds_pkt_valid = (demux_select== 9'd15) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress16_ds_pkt_valid = (demux_select== 9'd16) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress17_ds_pkt_valid = (demux_select== 9'd17) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress18_ds_pkt_valid = (demux_select== 9'd18) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress19_ds_pkt_valid = (demux_select== 9'd19) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress20_ds_pkt_valid = (demux_select== 9'd20) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress21_ds_pkt_valid = (demux_select== 9'd21) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress22_ds_pkt_valid = (demux_select== 9'd22) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress23_ds_pkt_valid = (demux_select== 9'd23) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress24_ds_pkt_valid = (demux_select== 9'd24) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress25_ds_pkt_valid = (demux_select== 9'd25) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress26_ds_pkt_valid = (demux_select== 9'd26) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress27_ds_pkt_valid = (demux_select== 9'd27) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress28_ds_pkt_valid = (demux_select== 9'd28) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress29_ds_pkt_valid = (demux_select== 9'd29) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress30_ds_pkt_valid = (demux_select== 9'd30) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress31_ds_pkt_valid = (demux_select== 9'd31) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress32_ds_pkt_valid = (demux_select== 9'd32) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress33_ds_pkt_valid = (demux_select== 9'd33) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress34_ds_pkt_valid = (demux_select== 9'd34) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress35_ds_pkt_valid = (demux_select== 9'd35) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress36_ds_pkt_valid = (demux_select== 9'd36) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress37_ds_pkt_valid = (demux_select== 9'd37) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress38_ds_pkt_valid = (demux_select== 9'd38) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress39_ds_pkt_valid = (demux_select== 9'd39) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress40_ds_pkt_valid = (demux_select== 9'd40) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress41_ds_pkt_valid = (demux_select== 9'd41) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress42_ds_pkt_valid = (demux_select== 9'd42) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress43_ds_pkt_valid = (demux_select== 9'd43) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress44_ds_pkt_valid = (demux_select== 9'd44) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress45_ds_pkt_valid = (demux_select== 9'd45) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress46_ds_pkt_valid = (demux_select== 9'd46) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress47_ds_pkt_valid = (demux_select== 9'd47) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress48_ds_pkt_valid = (demux_select== 9'd48) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress49_ds_pkt_valid = (demux_select== 9'd49) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress50_ds_pkt_valid = (demux_select== 9'd50) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress51_ds_pkt_valid = (demux_select== 9'd51) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress52_ds_pkt_valid = (demux_select== 9'd52) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress53_ds_pkt_valid = (demux_select== 9'd53) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress54_ds_pkt_valid = (demux_select== 9'd54) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress55_ds_pkt_valid = (demux_select== 9'd55) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress56_ds_pkt_valid = (demux_select== 9'd56) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress57_ds_pkt_valid = (demux_select== 9'd57) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress58_ds_pkt_valid = (demux_select== 9'd58) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress59_ds_pkt_valid = (demux_select== 9'd59) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress60_ds_pkt_valid = (demux_select== 9'd60) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress61_ds_pkt_valid = (demux_select== 9'd61) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress62_ds_pkt_valid = (demux_select== 9'd62) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress63_ds_pkt_valid = (demux_select== 9'd63) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress64_ds_pkt_valid = (demux_select== 9'd64) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress65_ds_pkt_valid = (demux_select== 9'd65) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress66_ds_pkt_valid = (demux_select== 9'd66) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress67_ds_pkt_valid = (demux_select== 9'd67) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress68_ds_pkt_valid = (demux_select== 9'd68) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress69_ds_pkt_valid = (demux_select== 9'd69) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress70_ds_pkt_valid = (demux_select== 9'd70) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress71_ds_pkt_valid = (demux_select== 9'd71) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress72_ds_pkt_valid = (demux_select== 9'd72) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress73_ds_pkt_valid = (demux_select== 9'd73) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress74_ds_pkt_valid = (demux_select== 9'd74) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress75_ds_pkt_valid = (demux_select== 9'd75) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress76_ds_pkt_valid = (demux_select== 9'd76) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress77_ds_pkt_valid = (demux_select== 9'd77) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress78_ds_pkt_valid = (demux_select== 9'd78) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress79_ds_pkt_valid = (demux_select== 9'd79) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress80_ds_pkt_valid = (demux_select== 9'd80) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress81_ds_pkt_valid = (demux_select== 9'd81) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress82_ds_pkt_valid = (demux_select== 9'd82) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress83_ds_pkt_valid = (demux_select== 9'd83) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress84_ds_pkt_valid = (demux_select== 9'd84) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress85_ds_pkt_valid = (demux_select== 9'd85) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress86_ds_pkt_valid = (demux_select== 9'd86) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress87_ds_pkt_valid = (demux_select== 9'd87) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress88_ds_pkt_valid = (demux_select== 9'd88) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress89_ds_pkt_valid = (demux_select== 9'd89) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress90_ds_pkt_valid = (demux_select== 9'd90) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress91_ds_pkt_valid = (demux_select== 9'd91) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress92_ds_pkt_valid = (demux_select== 9'd92) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress93_ds_pkt_valid = (demux_select== 9'd93) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress94_ds_pkt_valid = (demux_select== 9'd94) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress95_ds_pkt_valid = (demux_select== 9'd95) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress96_ds_pkt_valid = (demux_select== 9'd96) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress97_ds_pkt_valid = (demux_select== 9'd97) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress98_ds_pkt_valid = (demux_select== 9'd98) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress99_ds_pkt_valid = (demux_select== 9'd99) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress100_ds_pkt_valid = (demux_select== 9'd100) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress101_ds_pkt_valid = (demux_select== 9'd101) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress102_ds_pkt_valid = (demux_select== 9'd102) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress103_ds_pkt_valid = (demux_select== 9'd103) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress104_ds_pkt_valid = (demux_select== 9'd104) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress105_ds_pkt_valid = (demux_select== 9'd105) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress106_ds_pkt_valid = (demux_select== 9'd106) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress107_ds_pkt_valid = (demux_select== 9'd107) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress108_ds_pkt_valid = (demux_select== 9'd108) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress109_ds_pkt_valid = (demux_select== 9'd109) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress110_ds_pkt_valid = (demux_select== 9'd110) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress111_ds_pkt_valid = (demux_select== 9'd111) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress112_ds_pkt_valid = (demux_select== 9'd112) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress113_ds_pkt_valid = (demux_select== 9'd113) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress114_ds_pkt_valid = (demux_select== 9'd114) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress115_ds_pkt_valid = (demux_select== 9'd115) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress116_ds_pkt_valid = (demux_select== 9'd116) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress117_ds_pkt_valid = (demux_select== 9'd117) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress118_ds_pkt_valid = (demux_select== 9'd118) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress119_ds_pkt_valid = (demux_select== 9'd119) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress120_ds_pkt_valid = (demux_select== 9'd120) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress121_ds_pkt_valid = (demux_select== 9'd121) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress122_ds_pkt_valid = (demux_select== 9'd122) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress123_ds_pkt_valid = (demux_select== 9'd123) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress124_ds_pkt_valid = (demux_select== 9'd124) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress125_ds_pkt_valid = (demux_select== 9'd125) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress126_ds_pkt_valid = (demux_select== 9'd126) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress127_ds_pkt_valid = (demux_select== 9'd127) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress128_ds_pkt_valid = (demux_select== 9'd128) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress129_ds_pkt_valid = (demux_select== 9'd129) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress130_ds_pkt_valid = (demux_select== 9'd130) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress131_ds_pkt_valid = (demux_select== 9'd131) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress132_ds_pkt_valid = (demux_select== 9'd132) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress133_ds_pkt_valid = (demux_select== 9'd133) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress134_ds_pkt_valid = (demux_select== 9'd134) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress135_ds_pkt_valid = (demux_select== 9'd135) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress136_ds_pkt_valid = (demux_select== 9'd136) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress137_ds_pkt_valid = (demux_select== 9'd137) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress138_ds_pkt_valid = (demux_select== 9'd138) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress139_ds_pkt_valid = (demux_select== 9'd139) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress140_ds_pkt_valid = (demux_select== 9'd140) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress141_ds_pkt_valid = (demux_select== 9'd141) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress142_ds_pkt_valid = (demux_select== 9'd142) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress143_ds_pkt_valid = (demux_select== 9'd143) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress144_ds_pkt_valid = (demux_select== 9'd144) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress145_ds_pkt_valid = (demux_select== 9'd145) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress146_ds_pkt_valid = (demux_select== 9'd146) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress147_ds_pkt_valid = (demux_select== 9'd147) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress148_ds_pkt_valid = (demux_select== 9'd148) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress149_ds_pkt_valid = (demux_select== 9'd149) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress150_ds_pkt_valid = (demux_select== 9'd150) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress151_ds_pkt_valid = (demux_select== 9'd151) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress152_ds_pkt_valid = (demux_select== 9'd152) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress153_ds_pkt_valid = (demux_select== 9'd153) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress154_ds_pkt_valid = (demux_select== 9'd154) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress155_ds_pkt_valid = (demux_select== 9'd155) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress156_ds_pkt_valid = (demux_select== 9'd156) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress157_ds_pkt_valid = (demux_select== 9'd157) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress158_ds_pkt_valid = (demux_select== 9'd158) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress159_ds_pkt_valid = (demux_select== 9'd159) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress160_ds_pkt_valid = (demux_select== 9'd160) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress161_ds_pkt_valid = (demux_select== 9'd161) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress162_ds_pkt_valid = (demux_select== 9'd162) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress163_ds_pkt_valid = (demux_select== 9'd163) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress164_ds_pkt_valid = (demux_select== 9'd164) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress165_ds_pkt_valid = (demux_select== 9'd165) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress166_ds_pkt_valid = (demux_select== 9'd166) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress167_ds_pkt_valid = (demux_select== 9'd167) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress168_ds_pkt_valid = (demux_select== 9'd168) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress169_ds_pkt_valid = (demux_select== 9'd169) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress170_ds_pkt_valid = (demux_select== 9'd170) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress171_ds_pkt_valid = (demux_select== 9'd171) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress172_ds_pkt_valid = (demux_select== 9'd172) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress173_ds_pkt_valid = (demux_select== 9'd173) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress174_ds_pkt_valid = (demux_select== 9'd174) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress175_ds_pkt_valid = (demux_select== 9'd175) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress176_ds_pkt_valid = (demux_select== 9'd176) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress177_ds_pkt_valid = (demux_select== 9'd177) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress178_ds_pkt_valid = (demux_select== 9'd178) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress179_ds_pkt_valid = (demux_select== 9'd179) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress180_ds_pkt_valid = (demux_select== 9'd180) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress181_ds_pkt_valid = (demux_select== 9'd181) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress182_ds_pkt_valid = (demux_select== 9'd182) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress183_ds_pkt_valid = (demux_select== 9'd183) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress184_ds_pkt_valid = (demux_select== 9'd184) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress185_ds_pkt_valid = (demux_select== 9'd185) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress186_ds_pkt_valid = (demux_select== 9'd186) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress187_ds_pkt_valid = (demux_select== 9'd187) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress188_ds_pkt_valid = (demux_select== 9'd188) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress189_ds_pkt_valid = (demux_select== 9'd189) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress190_ds_pkt_valid = (demux_select== 9'd190) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress191_ds_pkt_valid = (demux_select== 9'd191) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress192_ds_pkt_valid = (demux_select== 9'd192) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress193_ds_pkt_valid = (demux_select== 9'd193) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress194_ds_pkt_valid = (demux_select== 9'd194) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress195_ds_pkt_valid = (demux_select== 9'd195) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress196_ds_pkt_valid = (demux_select== 9'd196) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress197_ds_pkt_valid = (demux_select== 9'd197) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress198_ds_pkt_valid = (demux_select== 9'd198) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress199_ds_pkt_valid = (demux_select== 9'd199) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress200_ds_pkt_valid = (demux_select== 9'd200) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress201_ds_pkt_valid = (demux_select== 9'd201) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress202_ds_pkt_valid = (demux_select== 9'd202) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress203_ds_pkt_valid = (demux_select== 9'd203) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress204_ds_pkt_valid = (demux_select== 9'd204) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress205_ds_pkt_valid = (demux_select== 9'd205) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress206_ds_pkt_valid = (demux_select== 9'd206) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress207_ds_pkt_valid = (demux_select== 9'd207) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress208_ds_pkt_valid = (demux_select== 9'd208) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress209_ds_pkt_valid = (demux_select== 9'd209) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress210_ds_pkt_valid = (demux_select== 9'd210) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress211_ds_pkt_valid = (demux_select== 9'd211) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress212_ds_pkt_valid = (demux_select== 9'd212) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress213_ds_pkt_valid = (demux_select== 9'd213) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress214_ds_pkt_valid = (demux_select== 9'd214) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress215_ds_pkt_valid = (demux_select== 9'd215) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress216_ds_pkt_valid = (demux_select== 9'd216) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress217_ds_pkt_valid = (demux_select== 9'd217) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress218_ds_pkt_valid = (demux_select== 9'd218) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress219_ds_pkt_valid = (demux_select== 9'd219) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress220_ds_pkt_valid = (demux_select== 9'd220) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress221_ds_pkt_valid = (demux_select== 9'd221) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress222_ds_pkt_valid = (demux_select== 9'd222) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress223_ds_pkt_valid = (demux_select== 9'd223) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress224_ds_pkt_valid = (demux_select== 9'd224) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress225_ds_pkt_valid = (demux_select== 9'd225) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress226_ds_pkt_valid = (demux_select== 9'd226) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress227_ds_pkt_valid = (demux_select== 9'd227) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress228_ds_pkt_valid = (demux_select== 9'd228) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress229_ds_pkt_valid = (demux_select== 9'd229) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress230_ds_pkt_valid = (demux_select== 9'd230) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress231_ds_pkt_valid = (demux_select== 9'd231) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress232_ds_pkt_valid = (demux_select== 9'd232) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress233_ds_pkt_valid = (demux_select== 9'd233) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress234_ds_pkt_valid = (demux_select== 9'd234) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress235_ds_pkt_valid = (demux_select== 9'd235) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress236_ds_pkt_valid = (demux_select== 9'd236) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress237_ds_pkt_valid = (demux_select== 9'd237) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress238_ds_pkt_valid = (demux_select== 9'd238) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress239_ds_pkt_valid = (demux_select== 9'd239) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress240_ds_pkt_valid = (demux_select== 9'd240) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress241_ds_pkt_valid = (demux_select== 9'd241) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress242_ds_pkt_valid = (demux_select== 9'd242) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress243_ds_pkt_valid = (demux_select== 9'd243) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress244_ds_pkt_valid = (demux_select== 9'd244) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress245_ds_pkt_valid = (demux_select== 9'd245) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress246_ds_pkt_valid = (demux_select== 9'd246) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress247_ds_pkt_valid = (demux_select== 9'd247) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress248_ds_pkt_valid = (demux_select== 9'd248) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress249_ds_pkt_valid = (demux_select== 9'd249) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress250_ds_pkt_valid = (demux_select== 9'd250) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress251_ds_pkt_valid = (demux_select== 9'd251) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress252_ds_pkt_valid = (demux_select== 9'd252) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress253_ds_pkt_valid = (demux_select== 9'd253) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress254_ds_pkt_valid = (demux_select== 9'd254) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress255_ds_pkt_valid = (demux_select== 9'd255) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress256_ds_pkt_valid = (demux_select== 9'd256) ? ingress_ds_pkt_valid : 9'd0;
wire assign egress257_ds_pkt_valid = (demux_select== 9'd257) ? ingress_ds_pkt_valid : 9'd0;

wire assign ingress_ds_pkt_ready          =
                                           ((demux_select== 9'd0) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd1) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd2) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd3) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd4) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd5) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd6) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd7) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd8) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd9) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd10) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd11) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd12) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd13) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd14) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd15) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd16) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd17) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd18) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd19) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd20) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd21) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd22) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd23) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd24) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd25) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd26) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd27) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd28) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd29) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd30) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd31) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd32) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd33) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd34) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd35) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd36) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd37) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd38) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd39) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd40) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd41) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd42) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd43) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd44) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd45) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd46) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd47) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd48) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd49) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd50) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd51) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd52) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd53) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd54) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd55) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd56) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd57) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd58) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd59) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd60) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd61) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd62) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd63) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd64) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd65) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd66) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd67) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd68) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd69) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd70) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd71) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd72) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd73) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd74) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd75) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd76) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd77) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd78) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd79) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd80) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd81) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd82) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd83) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd84) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd85) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd86) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd87) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd88) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd89) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd90) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd91) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd92) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd93) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd94) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd95) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd96) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd97) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd98) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd99) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd100) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd101) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd102) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd103) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd104) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd105) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd106) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd107) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd108) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd109) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd110) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd111) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd112) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd113) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd114) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd115) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd116) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd117) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd118) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd119) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd120) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd121) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd122) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd123) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd124) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd125) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd126) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd127) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd128) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd129) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd130) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd131) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd132) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd133) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd134) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd135) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd136) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd137) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd138) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd139) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd140) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd141) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd142) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd143) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd144) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd145) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd146) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd147) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd148) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd149) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd150) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd151) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd152) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd153) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd154) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd155) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd156) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd157) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd158) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd159) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd160) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd161) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd162) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd163) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd164) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd165) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd166) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd167) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd168) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd169) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd170) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd171) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd172) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd173) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd174) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd175) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd176) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd177) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd178) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd179) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd180) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd181) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd182) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd183) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd184) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd185) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd186) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd187) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd188) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd189) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd190) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd191) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd192) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd193) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd194) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd195) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd196) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd197) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd198) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd199) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd200) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd201) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd202) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd203) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd204) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd205) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd206) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd207) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd208) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd209) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd210) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd211) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd212) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd213) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd214) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd215) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd216) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd217) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd218) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd219) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd220) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd221) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd222) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd223) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd224) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd225) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd226) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd227) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd228) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd229) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd230) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd231) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd232) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd233) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd234) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd235) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd236) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd237) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd238) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd239) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd240) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd241) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd242) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd243) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd244) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd245) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd246) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd247) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd248) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd249) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd250) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd251) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd252) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd253) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd254) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd255) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd256) ? egress1_ds_pkt_ready ? 1'b0) | 
                                           ((demux_select== 9'd257) ? egress1_ds_pkt_ready ? 1'b0) | 
                                            1'b0;



endmodule
