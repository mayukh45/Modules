
module AH_CAM_1100_20_15 (wdata
,wvalid
,wready
,sdata
,svalid
,smatch
,sin);

input [19:0] wdata;
input wvalid;
output wready;
input [19:0] sdata;
input svalid;
input smatch;
input [14:0] sin;

wire [10:0] internal_wr_ptr;
req  [11:0] wr_loc_counter;
        req  [19:0] cam_loc0;
req  [19:0] cam_loc1;
req  [19:0] cam_loc2;
req  [19:0] cam_loc3;
req  [19:0] cam_loc4;
req  [19:0] cam_loc5;
req  [19:0] cam_loc6;
req  [19:0] cam_loc7;
req  [19:0] cam_loc8;
req  [19:0] cam_loc9;
req  [19:0] cam_loc10;
req  [19:0] cam_loc11;
req  [19:0] cam_loc12;
req  [19:0] cam_loc13;
req  [19:0] cam_loc14;
req  [19:0] cam_loc15;
req  [19:0] cam_loc16;
req  [19:0] cam_loc17;
req  [19:0] cam_loc18;
req  [19:0] cam_loc19;
req  [19:0] cam_loc20;
req  [19:0] cam_loc21;
req  [19:0] cam_loc22;
req  [19:0] cam_loc23;
req  [19:0] cam_loc24;
req  [19:0] cam_loc25;
req  [19:0] cam_loc26;
req  [19:0] cam_loc27;
req  [19:0] cam_loc28;
req  [19:0] cam_loc29;
req  [19:0] cam_loc30;
req  [19:0] cam_loc31;
req  [19:0] cam_loc32;
req  [19:0] cam_loc33;
req  [19:0] cam_loc34;
req  [19:0] cam_loc35;
req  [19:0] cam_loc36;
req  [19:0] cam_loc37;
req  [19:0] cam_loc38;
req  [19:0] cam_loc39;
req  [19:0] cam_loc40;
req  [19:0] cam_loc41;
req  [19:0] cam_loc42;
req  [19:0] cam_loc43;
req  [19:0] cam_loc44;
req  [19:0] cam_loc45;
req  [19:0] cam_loc46;
req  [19:0] cam_loc47;
req  [19:0] cam_loc48;
req  [19:0] cam_loc49;
req  [19:0] cam_loc50;
req  [19:0] cam_loc51;
req  [19:0] cam_loc52;
req  [19:0] cam_loc53;
req  [19:0] cam_loc54;
req  [19:0] cam_loc55;
req  [19:0] cam_loc56;
req  [19:0] cam_loc57;
req  [19:0] cam_loc58;
req  [19:0] cam_loc59;
req  [19:0] cam_loc60;
req  [19:0] cam_loc61;
req  [19:0] cam_loc62;
req  [19:0] cam_loc63;
req  [19:0] cam_loc64;
req  [19:0] cam_loc65;
req  [19:0] cam_loc66;
req  [19:0] cam_loc67;
req  [19:0] cam_loc68;
req  [19:0] cam_loc69;
req  [19:0] cam_loc70;
req  [19:0] cam_loc71;
req  [19:0] cam_loc72;
req  [19:0] cam_loc73;
req  [19:0] cam_loc74;
req  [19:0] cam_loc75;
req  [19:0] cam_loc76;
req  [19:0] cam_loc77;
req  [19:0] cam_loc78;
req  [19:0] cam_loc79;
req  [19:0] cam_loc80;
req  [19:0] cam_loc81;
req  [19:0] cam_loc82;
req  [19:0] cam_loc83;
req  [19:0] cam_loc84;
req  [19:0] cam_loc85;
req  [19:0] cam_loc86;
req  [19:0] cam_loc87;
req  [19:0] cam_loc88;
req  [19:0] cam_loc89;
req  [19:0] cam_loc90;
req  [19:0] cam_loc91;
req  [19:0] cam_loc92;
req  [19:0] cam_loc93;
req  [19:0] cam_loc94;
req  [19:0] cam_loc95;
req  [19:0] cam_loc96;
req  [19:0] cam_loc97;
req  [19:0] cam_loc98;
req  [19:0] cam_loc99;
req  [19:0] cam_loc100;
req  [19:0] cam_loc101;
req  [19:0] cam_loc102;
req  [19:0] cam_loc103;
req  [19:0] cam_loc104;
req  [19:0] cam_loc105;
req  [19:0] cam_loc106;
req  [19:0] cam_loc107;
req  [19:0] cam_loc108;
req  [19:0] cam_loc109;
req  [19:0] cam_loc110;
req  [19:0] cam_loc111;
req  [19:0] cam_loc112;
req  [19:0] cam_loc113;
req  [19:0] cam_loc114;
req  [19:0] cam_loc115;
req  [19:0] cam_loc116;
req  [19:0] cam_loc117;
req  [19:0] cam_loc118;
req  [19:0] cam_loc119;
req  [19:0] cam_loc120;
req  [19:0] cam_loc121;
req  [19:0] cam_loc122;
req  [19:0] cam_loc123;
req  [19:0] cam_loc124;
req  [19:0] cam_loc125;
req  [19:0] cam_loc126;
req  [19:0] cam_loc127;
req  [19:0] cam_loc128;
req  [19:0] cam_loc129;
req  [19:0] cam_loc130;
req  [19:0] cam_loc131;
req  [19:0] cam_loc132;
req  [19:0] cam_loc133;
req  [19:0] cam_loc134;
req  [19:0] cam_loc135;
req  [19:0] cam_loc136;
req  [19:0] cam_loc137;
req  [19:0] cam_loc138;
req  [19:0] cam_loc139;
req  [19:0] cam_loc140;
req  [19:0] cam_loc141;
req  [19:0] cam_loc142;
req  [19:0] cam_loc143;
req  [19:0] cam_loc144;
req  [19:0] cam_loc145;
req  [19:0] cam_loc146;
req  [19:0] cam_loc147;
req  [19:0] cam_loc148;
req  [19:0] cam_loc149;
req  [19:0] cam_loc150;
req  [19:0] cam_loc151;
req  [19:0] cam_loc152;
req  [19:0] cam_loc153;
req  [19:0] cam_loc154;
req  [19:0] cam_loc155;
req  [19:0] cam_loc156;
req  [19:0] cam_loc157;
req  [19:0] cam_loc158;
req  [19:0] cam_loc159;
req  [19:0] cam_loc160;
req  [19:0] cam_loc161;
req  [19:0] cam_loc162;
req  [19:0] cam_loc163;
req  [19:0] cam_loc164;
req  [19:0] cam_loc165;
req  [19:0] cam_loc166;
req  [19:0] cam_loc167;
req  [19:0] cam_loc168;
req  [19:0] cam_loc169;
req  [19:0] cam_loc170;
req  [19:0] cam_loc171;
req  [19:0] cam_loc172;
req  [19:0] cam_loc173;
req  [19:0] cam_loc174;
req  [19:0] cam_loc175;
req  [19:0] cam_loc176;
req  [19:0] cam_loc177;
req  [19:0] cam_loc178;
req  [19:0] cam_loc179;
req  [19:0] cam_loc180;
req  [19:0] cam_loc181;
req  [19:0] cam_loc182;
req  [19:0] cam_loc183;
req  [19:0] cam_loc184;
req  [19:0] cam_loc185;
req  [19:0] cam_loc186;
req  [19:0] cam_loc187;
req  [19:0] cam_loc188;
req  [19:0] cam_loc189;
req  [19:0] cam_loc190;
req  [19:0] cam_loc191;
req  [19:0] cam_loc192;
req  [19:0] cam_loc193;
req  [19:0] cam_loc194;
req  [19:0] cam_loc195;
req  [19:0] cam_loc196;
req  [19:0] cam_loc197;
req  [19:0] cam_loc198;
req  [19:0] cam_loc199;
req  [19:0] cam_loc200;
req  [19:0] cam_loc201;
req  [19:0] cam_loc202;
req  [19:0] cam_loc203;
req  [19:0] cam_loc204;
req  [19:0] cam_loc205;
req  [19:0] cam_loc206;
req  [19:0] cam_loc207;
req  [19:0] cam_loc208;
req  [19:0] cam_loc209;
req  [19:0] cam_loc210;
req  [19:0] cam_loc211;
req  [19:0] cam_loc212;
req  [19:0] cam_loc213;
req  [19:0] cam_loc214;
req  [19:0] cam_loc215;
req  [19:0] cam_loc216;
req  [19:0] cam_loc217;
req  [19:0] cam_loc218;
req  [19:0] cam_loc219;
req  [19:0] cam_loc220;
req  [19:0] cam_loc221;
req  [19:0] cam_loc222;
req  [19:0] cam_loc223;
req  [19:0] cam_loc224;
req  [19:0] cam_loc225;
req  [19:0] cam_loc226;
req  [19:0] cam_loc227;
req  [19:0] cam_loc228;
req  [19:0] cam_loc229;
req  [19:0] cam_loc230;
req  [19:0] cam_loc231;
req  [19:0] cam_loc232;
req  [19:0] cam_loc233;
req  [19:0] cam_loc234;
req  [19:0] cam_loc235;
req  [19:0] cam_loc236;
req  [19:0] cam_loc237;
req  [19:0] cam_loc238;
req  [19:0] cam_loc239;
req  [19:0] cam_loc240;
req  [19:0] cam_loc241;
req  [19:0] cam_loc242;
req  [19:0] cam_loc243;
req  [19:0] cam_loc244;
req  [19:0] cam_loc245;
req  [19:0] cam_loc246;
req  [19:0] cam_loc247;
req  [19:0] cam_loc248;
req  [19:0] cam_loc249;
req  [19:0] cam_loc250;
req  [19:0] cam_loc251;
req  [19:0] cam_loc252;
req  [19:0] cam_loc253;
req  [19:0] cam_loc254;
req  [19:0] cam_loc255;
req  [19:0] cam_loc256;
req  [19:0] cam_loc257;
req  [19:0] cam_loc258;
req  [19:0] cam_loc259;
req  [19:0] cam_loc260;
req  [19:0] cam_loc261;
req  [19:0] cam_loc262;
req  [19:0] cam_loc263;
req  [19:0] cam_loc264;
req  [19:0] cam_loc265;
req  [19:0] cam_loc266;
req  [19:0] cam_loc267;
req  [19:0] cam_loc268;
req  [19:0] cam_loc269;
req  [19:0] cam_loc270;
req  [19:0] cam_loc271;
req  [19:0] cam_loc272;
req  [19:0] cam_loc273;
req  [19:0] cam_loc274;
req  [19:0] cam_loc275;
req  [19:0] cam_loc276;
req  [19:0] cam_loc277;
req  [19:0] cam_loc278;
req  [19:0] cam_loc279;
req  [19:0] cam_loc280;
req  [19:0] cam_loc281;
req  [19:0] cam_loc282;
req  [19:0] cam_loc283;
req  [19:0] cam_loc284;
req  [19:0] cam_loc285;
req  [19:0] cam_loc286;
req  [19:0] cam_loc287;
req  [19:0] cam_loc288;
req  [19:0] cam_loc289;
req  [19:0] cam_loc290;
req  [19:0] cam_loc291;
req  [19:0] cam_loc292;
req  [19:0] cam_loc293;
req  [19:0] cam_loc294;
req  [19:0] cam_loc295;
req  [19:0] cam_loc296;
req  [19:0] cam_loc297;
req  [19:0] cam_loc298;
req  [19:0] cam_loc299;
req  [19:0] cam_loc300;
req  [19:0] cam_loc301;
req  [19:0] cam_loc302;
req  [19:0] cam_loc303;
req  [19:0] cam_loc304;
req  [19:0] cam_loc305;
req  [19:0] cam_loc306;
req  [19:0] cam_loc307;
req  [19:0] cam_loc308;
req  [19:0] cam_loc309;
req  [19:0] cam_loc310;
req  [19:0] cam_loc311;
req  [19:0] cam_loc312;
req  [19:0] cam_loc313;
req  [19:0] cam_loc314;
req  [19:0] cam_loc315;
req  [19:0] cam_loc316;
req  [19:0] cam_loc317;
req  [19:0] cam_loc318;
req  [19:0] cam_loc319;
req  [19:0] cam_loc320;
req  [19:0] cam_loc321;
req  [19:0] cam_loc322;
req  [19:0] cam_loc323;
req  [19:0] cam_loc324;
req  [19:0] cam_loc325;
req  [19:0] cam_loc326;
req  [19:0] cam_loc327;
req  [19:0] cam_loc328;
req  [19:0] cam_loc329;
req  [19:0] cam_loc330;
req  [19:0] cam_loc331;
req  [19:0] cam_loc332;
req  [19:0] cam_loc333;
req  [19:0] cam_loc334;
req  [19:0] cam_loc335;
req  [19:0] cam_loc336;
req  [19:0] cam_loc337;
req  [19:0] cam_loc338;
req  [19:0] cam_loc339;
req  [19:0] cam_loc340;
req  [19:0] cam_loc341;
req  [19:0] cam_loc342;
req  [19:0] cam_loc343;
req  [19:0] cam_loc344;
req  [19:0] cam_loc345;
req  [19:0] cam_loc346;
req  [19:0] cam_loc347;
req  [19:0] cam_loc348;
req  [19:0] cam_loc349;
req  [19:0] cam_loc350;
req  [19:0] cam_loc351;
req  [19:0] cam_loc352;
req  [19:0] cam_loc353;
req  [19:0] cam_loc354;
req  [19:0] cam_loc355;
req  [19:0] cam_loc356;
req  [19:0] cam_loc357;
req  [19:0] cam_loc358;
req  [19:0] cam_loc359;
req  [19:0] cam_loc360;
req  [19:0] cam_loc361;
req  [19:0] cam_loc362;
req  [19:0] cam_loc363;
req  [19:0] cam_loc364;
req  [19:0] cam_loc365;
req  [19:0] cam_loc366;
req  [19:0] cam_loc367;
req  [19:0] cam_loc368;
req  [19:0] cam_loc369;
req  [19:0] cam_loc370;
req  [19:0] cam_loc371;
req  [19:0] cam_loc372;
req  [19:0] cam_loc373;
req  [19:0] cam_loc374;
req  [19:0] cam_loc375;
req  [19:0] cam_loc376;
req  [19:0] cam_loc377;
req  [19:0] cam_loc378;
req  [19:0] cam_loc379;
req  [19:0] cam_loc380;
req  [19:0] cam_loc381;
req  [19:0] cam_loc382;
req  [19:0] cam_loc383;
req  [19:0] cam_loc384;
req  [19:0] cam_loc385;
req  [19:0] cam_loc386;
req  [19:0] cam_loc387;
req  [19:0] cam_loc388;
req  [19:0] cam_loc389;
req  [19:0] cam_loc390;
req  [19:0] cam_loc391;
req  [19:0] cam_loc392;
req  [19:0] cam_loc393;
req  [19:0] cam_loc394;
req  [19:0] cam_loc395;
req  [19:0] cam_loc396;
req  [19:0] cam_loc397;
req  [19:0] cam_loc398;
req  [19:0] cam_loc399;
req  [19:0] cam_loc400;
req  [19:0] cam_loc401;
req  [19:0] cam_loc402;
req  [19:0] cam_loc403;
req  [19:0] cam_loc404;
req  [19:0] cam_loc405;
req  [19:0] cam_loc406;
req  [19:0] cam_loc407;
req  [19:0] cam_loc408;
req  [19:0] cam_loc409;
req  [19:0] cam_loc410;
req  [19:0] cam_loc411;
req  [19:0] cam_loc412;
req  [19:0] cam_loc413;
req  [19:0] cam_loc414;
req  [19:0] cam_loc415;
req  [19:0] cam_loc416;
req  [19:0] cam_loc417;
req  [19:0] cam_loc418;
req  [19:0] cam_loc419;
req  [19:0] cam_loc420;
req  [19:0] cam_loc421;
req  [19:0] cam_loc422;
req  [19:0] cam_loc423;
req  [19:0] cam_loc424;
req  [19:0] cam_loc425;
req  [19:0] cam_loc426;
req  [19:0] cam_loc427;
req  [19:0] cam_loc428;
req  [19:0] cam_loc429;
req  [19:0] cam_loc430;
req  [19:0] cam_loc431;
req  [19:0] cam_loc432;
req  [19:0] cam_loc433;
req  [19:0] cam_loc434;
req  [19:0] cam_loc435;
req  [19:0] cam_loc436;
req  [19:0] cam_loc437;
req  [19:0] cam_loc438;
req  [19:0] cam_loc439;
req  [19:0] cam_loc440;
req  [19:0] cam_loc441;
req  [19:0] cam_loc442;
req  [19:0] cam_loc443;
req  [19:0] cam_loc444;
req  [19:0] cam_loc445;
req  [19:0] cam_loc446;
req  [19:0] cam_loc447;
req  [19:0] cam_loc448;
req  [19:0] cam_loc449;
req  [19:0] cam_loc450;
req  [19:0] cam_loc451;
req  [19:0] cam_loc452;
req  [19:0] cam_loc453;
req  [19:0] cam_loc454;
req  [19:0] cam_loc455;
req  [19:0] cam_loc456;
req  [19:0] cam_loc457;
req  [19:0] cam_loc458;
req  [19:0] cam_loc459;
req  [19:0] cam_loc460;
req  [19:0] cam_loc461;
req  [19:0] cam_loc462;
req  [19:0] cam_loc463;
req  [19:0] cam_loc464;
req  [19:0] cam_loc465;
req  [19:0] cam_loc466;
req  [19:0] cam_loc467;
req  [19:0] cam_loc468;
req  [19:0] cam_loc469;
req  [19:0] cam_loc470;
req  [19:0] cam_loc471;
req  [19:0] cam_loc472;
req  [19:0] cam_loc473;
req  [19:0] cam_loc474;
req  [19:0] cam_loc475;
req  [19:0] cam_loc476;
req  [19:0] cam_loc477;
req  [19:0] cam_loc478;
req  [19:0] cam_loc479;
req  [19:0] cam_loc480;
req  [19:0] cam_loc481;
req  [19:0] cam_loc482;
req  [19:0] cam_loc483;
req  [19:0] cam_loc484;
req  [19:0] cam_loc485;
req  [19:0] cam_loc486;
req  [19:0] cam_loc487;
req  [19:0] cam_loc488;
req  [19:0] cam_loc489;
req  [19:0] cam_loc490;
req  [19:0] cam_loc491;
req  [19:0] cam_loc492;
req  [19:0] cam_loc493;
req  [19:0] cam_loc494;
req  [19:0] cam_loc495;
req  [19:0] cam_loc496;
req  [19:0] cam_loc497;
req  [19:0] cam_loc498;
req  [19:0] cam_loc499;
req  [19:0] cam_loc500;
req  [19:0] cam_loc501;
req  [19:0] cam_loc502;
req  [19:0] cam_loc503;
req  [19:0] cam_loc504;
req  [19:0] cam_loc505;
req  [19:0] cam_loc506;
req  [19:0] cam_loc507;
req  [19:0] cam_loc508;
req  [19:0] cam_loc509;
req  [19:0] cam_loc510;
req  [19:0] cam_loc511;
req  [19:0] cam_loc512;
req  [19:0] cam_loc513;
req  [19:0] cam_loc514;
req  [19:0] cam_loc515;
req  [19:0] cam_loc516;
req  [19:0] cam_loc517;
req  [19:0] cam_loc518;
req  [19:0] cam_loc519;
req  [19:0] cam_loc520;
req  [19:0] cam_loc521;
req  [19:0] cam_loc522;
req  [19:0] cam_loc523;
req  [19:0] cam_loc524;
req  [19:0] cam_loc525;
req  [19:0] cam_loc526;
req  [19:0] cam_loc527;
req  [19:0] cam_loc528;
req  [19:0] cam_loc529;
req  [19:0] cam_loc530;
req  [19:0] cam_loc531;
req  [19:0] cam_loc532;
req  [19:0] cam_loc533;
req  [19:0] cam_loc534;
req  [19:0] cam_loc535;
req  [19:0] cam_loc536;
req  [19:0] cam_loc537;
req  [19:0] cam_loc538;
req  [19:0] cam_loc539;
req  [19:0] cam_loc540;
req  [19:0] cam_loc541;
req  [19:0] cam_loc542;
req  [19:0] cam_loc543;
req  [19:0] cam_loc544;
req  [19:0] cam_loc545;
req  [19:0] cam_loc546;
req  [19:0] cam_loc547;
req  [19:0] cam_loc548;
req  [19:0] cam_loc549;
req  [19:0] cam_loc550;
req  [19:0] cam_loc551;
req  [19:0] cam_loc552;
req  [19:0] cam_loc553;
req  [19:0] cam_loc554;
req  [19:0] cam_loc555;
req  [19:0] cam_loc556;
req  [19:0] cam_loc557;
req  [19:0] cam_loc558;
req  [19:0] cam_loc559;
req  [19:0] cam_loc560;
req  [19:0] cam_loc561;
req  [19:0] cam_loc562;
req  [19:0] cam_loc563;
req  [19:0] cam_loc564;
req  [19:0] cam_loc565;
req  [19:0] cam_loc566;
req  [19:0] cam_loc567;
req  [19:0] cam_loc568;
req  [19:0] cam_loc569;
req  [19:0] cam_loc570;
req  [19:0] cam_loc571;
req  [19:0] cam_loc572;
req  [19:0] cam_loc573;
req  [19:0] cam_loc574;
req  [19:0] cam_loc575;
req  [19:0] cam_loc576;
req  [19:0] cam_loc577;
req  [19:0] cam_loc578;
req  [19:0] cam_loc579;
req  [19:0] cam_loc580;
req  [19:0] cam_loc581;
req  [19:0] cam_loc582;
req  [19:0] cam_loc583;
req  [19:0] cam_loc584;
req  [19:0] cam_loc585;
req  [19:0] cam_loc586;
req  [19:0] cam_loc587;
req  [19:0] cam_loc588;
req  [19:0] cam_loc589;
req  [19:0] cam_loc590;
req  [19:0] cam_loc591;
req  [19:0] cam_loc592;
req  [19:0] cam_loc593;
req  [19:0] cam_loc594;
req  [19:0] cam_loc595;
req  [19:0] cam_loc596;
req  [19:0] cam_loc597;
req  [19:0] cam_loc598;
req  [19:0] cam_loc599;
req  [19:0] cam_loc600;
req  [19:0] cam_loc601;
req  [19:0] cam_loc602;
req  [19:0] cam_loc603;
req  [19:0] cam_loc604;
req  [19:0] cam_loc605;
req  [19:0] cam_loc606;
req  [19:0] cam_loc607;
req  [19:0] cam_loc608;
req  [19:0] cam_loc609;
req  [19:0] cam_loc610;
req  [19:0] cam_loc611;
req  [19:0] cam_loc612;
req  [19:0] cam_loc613;
req  [19:0] cam_loc614;
req  [19:0] cam_loc615;
req  [19:0] cam_loc616;
req  [19:0] cam_loc617;
req  [19:0] cam_loc618;
req  [19:0] cam_loc619;
req  [19:0] cam_loc620;
req  [19:0] cam_loc621;
req  [19:0] cam_loc622;
req  [19:0] cam_loc623;
req  [19:0] cam_loc624;
req  [19:0] cam_loc625;
req  [19:0] cam_loc626;
req  [19:0] cam_loc627;
req  [19:0] cam_loc628;
req  [19:0] cam_loc629;
req  [19:0] cam_loc630;
req  [19:0] cam_loc631;
req  [19:0] cam_loc632;
req  [19:0] cam_loc633;
req  [19:0] cam_loc634;
req  [19:0] cam_loc635;
req  [19:0] cam_loc636;
req  [19:0] cam_loc637;
req  [19:0] cam_loc638;
req  [19:0] cam_loc639;
req  [19:0] cam_loc640;
req  [19:0] cam_loc641;
req  [19:0] cam_loc642;
req  [19:0] cam_loc643;
req  [19:0] cam_loc644;
req  [19:0] cam_loc645;
req  [19:0] cam_loc646;
req  [19:0] cam_loc647;
req  [19:0] cam_loc648;
req  [19:0] cam_loc649;
req  [19:0] cam_loc650;
req  [19:0] cam_loc651;
req  [19:0] cam_loc652;
req  [19:0] cam_loc653;
req  [19:0] cam_loc654;
req  [19:0] cam_loc655;
req  [19:0] cam_loc656;
req  [19:0] cam_loc657;
req  [19:0] cam_loc658;
req  [19:0] cam_loc659;
req  [19:0] cam_loc660;
req  [19:0] cam_loc661;
req  [19:0] cam_loc662;
req  [19:0] cam_loc663;
req  [19:0] cam_loc664;
req  [19:0] cam_loc665;
req  [19:0] cam_loc666;
req  [19:0] cam_loc667;
req  [19:0] cam_loc668;
req  [19:0] cam_loc669;
req  [19:0] cam_loc670;
req  [19:0] cam_loc671;
req  [19:0] cam_loc672;
req  [19:0] cam_loc673;
req  [19:0] cam_loc674;
req  [19:0] cam_loc675;
req  [19:0] cam_loc676;
req  [19:0] cam_loc677;
req  [19:0] cam_loc678;
req  [19:0] cam_loc679;
req  [19:0] cam_loc680;
req  [19:0] cam_loc681;
req  [19:0] cam_loc682;
req  [19:0] cam_loc683;
req  [19:0] cam_loc684;
req  [19:0] cam_loc685;
req  [19:0] cam_loc686;
req  [19:0] cam_loc687;
req  [19:0] cam_loc688;
req  [19:0] cam_loc689;
req  [19:0] cam_loc690;
req  [19:0] cam_loc691;
req  [19:0] cam_loc692;
req  [19:0] cam_loc693;
req  [19:0] cam_loc694;
req  [19:0] cam_loc695;
req  [19:0] cam_loc696;
req  [19:0] cam_loc697;
req  [19:0] cam_loc698;
req  [19:0] cam_loc699;
req  [19:0] cam_loc700;
req  [19:0] cam_loc701;
req  [19:0] cam_loc702;
req  [19:0] cam_loc703;
req  [19:0] cam_loc704;
req  [19:0] cam_loc705;
req  [19:0] cam_loc706;
req  [19:0] cam_loc707;
req  [19:0] cam_loc708;
req  [19:0] cam_loc709;
req  [19:0] cam_loc710;
req  [19:0] cam_loc711;
req  [19:0] cam_loc712;
req  [19:0] cam_loc713;
req  [19:0] cam_loc714;
req  [19:0] cam_loc715;
req  [19:0] cam_loc716;
req  [19:0] cam_loc717;
req  [19:0] cam_loc718;
req  [19:0] cam_loc719;
req  [19:0] cam_loc720;
req  [19:0] cam_loc721;
req  [19:0] cam_loc722;
req  [19:0] cam_loc723;
req  [19:0] cam_loc724;
req  [19:0] cam_loc725;
req  [19:0] cam_loc726;
req  [19:0] cam_loc727;
req  [19:0] cam_loc728;
req  [19:0] cam_loc729;
req  [19:0] cam_loc730;
req  [19:0] cam_loc731;
req  [19:0] cam_loc732;
req  [19:0] cam_loc733;
req  [19:0] cam_loc734;
req  [19:0] cam_loc735;
req  [19:0] cam_loc736;
req  [19:0] cam_loc737;
req  [19:0] cam_loc738;
req  [19:0] cam_loc739;
req  [19:0] cam_loc740;
req  [19:0] cam_loc741;
req  [19:0] cam_loc742;
req  [19:0] cam_loc743;
req  [19:0] cam_loc744;
req  [19:0] cam_loc745;
req  [19:0] cam_loc746;
req  [19:0] cam_loc747;
req  [19:0] cam_loc748;
req  [19:0] cam_loc749;
req  [19:0] cam_loc750;
req  [19:0] cam_loc751;
req  [19:0] cam_loc752;
req  [19:0] cam_loc753;
req  [19:0] cam_loc754;
req  [19:0] cam_loc755;
req  [19:0] cam_loc756;
req  [19:0] cam_loc757;
req  [19:0] cam_loc758;
req  [19:0] cam_loc759;
req  [19:0] cam_loc760;
req  [19:0] cam_loc761;
req  [19:0] cam_loc762;
req  [19:0] cam_loc763;
req  [19:0] cam_loc764;
req  [19:0] cam_loc765;
req  [19:0] cam_loc766;
req  [19:0] cam_loc767;
req  [19:0] cam_loc768;
req  [19:0] cam_loc769;
req  [19:0] cam_loc770;
req  [19:0] cam_loc771;
req  [19:0] cam_loc772;
req  [19:0] cam_loc773;
req  [19:0] cam_loc774;
req  [19:0] cam_loc775;
req  [19:0] cam_loc776;
req  [19:0] cam_loc777;
req  [19:0] cam_loc778;
req  [19:0] cam_loc779;
req  [19:0] cam_loc780;
req  [19:0] cam_loc781;
req  [19:0] cam_loc782;
req  [19:0] cam_loc783;
req  [19:0] cam_loc784;
req  [19:0] cam_loc785;
req  [19:0] cam_loc786;
req  [19:0] cam_loc787;
req  [19:0] cam_loc788;
req  [19:0] cam_loc789;
req  [19:0] cam_loc790;
req  [19:0] cam_loc791;
req  [19:0] cam_loc792;
req  [19:0] cam_loc793;
req  [19:0] cam_loc794;
req  [19:0] cam_loc795;
req  [19:0] cam_loc796;
req  [19:0] cam_loc797;
req  [19:0] cam_loc798;
req  [19:0] cam_loc799;
req  [19:0] cam_loc800;
req  [19:0] cam_loc801;
req  [19:0] cam_loc802;
req  [19:0] cam_loc803;
req  [19:0] cam_loc804;
req  [19:0] cam_loc805;
req  [19:0] cam_loc806;
req  [19:0] cam_loc807;
req  [19:0] cam_loc808;
req  [19:0] cam_loc809;
req  [19:0] cam_loc810;
req  [19:0] cam_loc811;
req  [19:0] cam_loc812;
req  [19:0] cam_loc813;
req  [19:0] cam_loc814;
req  [19:0] cam_loc815;
req  [19:0] cam_loc816;
req  [19:0] cam_loc817;
req  [19:0] cam_loc818;
req  [19:0] cam_loc819;
req  [19:0] cam_loc820;
req  [19:0] cam_loc821;
req  [19:0] cam_loc822;
req  [19:0] cam_loc823;
req  [19:0] cam_loc824;
req  [19:0] cam_loc825;
req  [19:0] cam_loc826;
req  [19:0] cam_loc827;
req  [19:0] cam_loc828;
req  [19:0] cam_loc829;
req  [19:0] cam_loc830;
req  [19:0] cam_loc831;
req  [19:0] cam_loc832;
req  [19:0] cam_loc833;
req  [19:0] cam_loc834;
req  [19:0] cam_loc835;
req  [19:0] cam_loc836;
req  [19:0] cam_loc837;
req  [19:0] cam_loc838;
req  [19:0] cam_loc839;
req  [19:0] cam_loc840;
req  [19:0] cam_loc841;
req  [19:0] cam_loc842;
req  [19:0] cam_loc843;
req  [19:0] cam_loc844;
req  [19:0] cam_loc845;
req  [19:0] cam_loc846;
req  [19:0] cam_loc847;
req  [19:0] cam_loc848;
req  [19:0] cam_loc849;
req  [19:0] cam_loc850;
req  [19:0] cam_loc851;
req  [19:0] cam_loc852;
req  [19:0] cam_loc853;
req  [19:0] cam_loc854;
req  [19:0] cam_loc855;
req  [19:0] cam_loc856;
req  [19:0] cam_loc857;
req  [19:0] cam_loc858;
req  [19:0] cam_loc859;
req  [19:0] cam_loc860;
req  [19:0] cam_loc861;
req  [19:0] cam_loc862;
req  [19:0] cam_loc863;
req  [19:0] cam_loc864;
req  [19:0] cam_loc865;
req  [19:0] cam_loc866;
req  [19:0] cam_loc867;
req  [19:0] cam_loc868;
req  [19:0] cam_loc869;
req  [19:0] cam_loc870;
req  [19:0] cam_loc871;
req  [19:0] cam_loc872;
req  [19:0] cam_loc873;
req  [19:0] cam_loc874;
req  [19:0] cam_loc875;
req  [19:0] cam_loc876;
req  [19:0] cam_loc877;
req  [19:0] cam_loc878;
req  [19:0] cam_loc879;
req  [19:0] cam_loc880;
req  [19:0] cam_loc881;
req  [19:0] cam_loc882;
req  [19:0] cam_loc883;
req  [19:0] cam_loc884;
req  [19:0] cam_loc885;
req  [19:0] cam_loc886;
req  [19:0] cam_loc887;
req  [19:0] cam_loc888;
req  [19:0] cam_loc889;
req  [19:0] cam_loc890;
req  [19:0] cam_loc891;
req  [19:0] cam_loc892;
req  [19:0] cam_loc893;
req  [19:0] cam_loc894;
req  [19:0] cam_loc895;
req  [19:0] cam_loc896;
req  [19:0] cam_loc897;
req  [19:0] cam_loc898;
req  [19:0] cam_loc899;
req  [19:0] cam_loc900;
req  [19:0] cam_loc901;
req  [19:0] cam_loc902;
req  [19:0] cam_loc903;
req  [19:0] cam_loc904;
req  [19:0] cam_loc905;
req  [19:0] cam_loc906;
req  [19:0] cam_loc907;
req  [19:0] cam_loc908;
req  [19:0] cam_loc909;
req  [19:0] cam_loc910;
req  [19:0] cam_loc911;
req  [19:0] cam_loc912;
req  [19:0] cam_loc913;
req  [19:0] cam_loc914;
req  [19:0] cam_loc915;
req  [19:0] cam_loc916;
req  [19:0] cam_loc917;
req  [19:0] cam_loc918;
req  [19:0] cam_loc919;
req  [19:0] cam_loc920;
req  [19:0] cam_loc921;
req  [19:0] cam_loc922;
req  [19:0] cam_loc923;
req  [19:0] cam_loc924;
req  [19:0] cam_loc925;
req  [19:0] cam_loc926;
req  [19:0] cam_loc927;
req  [19:0] cam_loc928;
req  [19:0] cam_loc929;
req  [19:0] cam_loc930;
req  [19:0] cam_loc931;
req  [19:0] cam_loc932;
req  [19:0] cam_loc933;
req  [19:0] cam_loc934;
req  [19:0] cam_loc935;
req  [19:0] cam_loc936;
req  [19:0] cam_loc937;
req  [19:0] cam_loc938;
req  [19:0] cam_loc939;
req  [19:0] cam_loc940;
req  [19:0] cam_loc941;
req  [19:0] cam_loc942;
req  [19:0] cam_loc943;
req  [19:0] cam_loc944;
req  [19:0] cam_loc945;
req  [19:0] cam_loc946;
req  [19:0] cam_loc947;
req  [19:0] cam_loc948;
req  [19:0] cam_loc949;
req  [19:0] cam_loc950;
req  [19:0] cam_loc951;
req  [19:0] cam_loc952;
req  [19:0] cam_loc953;
req  [19:0] cam_loc954;
req  [19:0] cam_loc955;
req  [19:0] cam_loc956;
req  [19:0] cam_loc957;
req  [19:0] cam_loc958;
req  [19:0] cam_loc959;
req  [19:0] cam_loc960;
req  [19:0] cam_loc961;
req  [19:0] cam_loc962;
req  [19:0] cam_loc963;
req  [19:0] cam_loc964;
req  [19:0] cam_loc965;
req  [19:0] cam_loc966;
req  [19:0] cam_loc967;
req  [19:0] cam_loc968;
req  [19:0] cam_loc969;
req  [19:0] cam_loc970;
req  [19:0] cam_loc971;
req  [19:0] cam_loc972;
req  [19:0] cam_loc973;
req  [19:0] cam_loc974;
req  [19:0] cam_loc975;
req  [19:0] cam_loc976;
req  [19:0] cam_loc977;
req  [19:0] cam_loc978;
req  [19:0] cam_loc979;
req  [19:0] cam_loc980;
req  [19:0] cam_loc981;
req  [19:0] cam_loc982;
req  [19:0] cam_loc983;
req  [19:0] cam_loc984;
req  [19:0] cam_loc985;
req  [19:0] cam_loc986;
req  [19:0] cam_loc987;
req  [19:0] cam_loc988;
req  [19:0] cam_loc989;
req  [19:0] cam_loc990;
req  [19:0] cam_loc991;
req  [19:0] cam_loc992;
req  [19:0] cam_loc993;
req  [19:0] cam_loc994;
req  [19:0] cam_loc995;
req  [19:0] cam_loc996;
req  [19:0] cam_loc997;
req  [19:0] cam_loc998;
req  [19:0] cam_loc999;
req  [19:0] cam_loc1000;
req  [19:0] cam_loc1001;
req  [19:0] cam_loc1002;
req  [19:0] cam_loc1003;
req  [19:0] cam_loc1004;
req  [19:0] cam_loc1005;
req  [19:0] cam_loc1006;
req  [19:0] cam_loc1007;
req  [19:0] cam_loc1008;
req  [19:0] cam_loc1009;
req  [19:0] cam_loc1010;
req  [19:0] cam_loc1011;
req  [19:0] cam_loc1012;
req  [19:0] cam_loc1013;
req  [19:0] cam_loc1014;
req  [19:0] cam_loc1015;
req  [19:0] cam_loc1016;
req  [19:0] cam_loc1017;
req  [19:0] cam_loc1018;
req  [19:0] cam_loc1019;
req  [19:0] cam_loc1020;
req  [19:0] cam_loc1021;
req  [19:0] cam_loc1022;
req  [19:0] cam_loc1023;
req  [19:0] cam_loc1024;
req  [19:0] cam_loc1025;
req  [19:0] cam_loc1026;
req  [19:0] cam_loc1027;
req  [19:0] cam_loc1028;
req  [19:0] cam_loc1029;
req  [19:0] cam_loc1030;
req  [19:0] cam_loc1031;
req  [19:0] cam_loc1032;
req  [19:0] cam_loc1033;
req  [19:0] cam_loc1034;
req  [19:0] cam_loc1035;
req  [19:0] cam_loc1036;
req  [19:0] cam_loc1037;
req  [19:0] cam_loc1038;
req  [19:0] cam_loc1039;
req  [19:0] cam_loc1040;
req  [19:0] cam_loc1041;
req  [19:0] cam_loc1042;
req  [19:0] cam_loc1043;
req  [19:0] cam_loc1044;
req  [19:0] cam_loc1045;
req  [19:0] cam_loc1046;
req  [19:0] cam_loc1047;
req  [19:0] cam_loc1048;
req  [19:0] cam_loc1049;
req  [19:0] cam_loc1050;
req  [19:0] cam_loc1051;
req  [19:0] cam_loc1052;
req  [19:0] cam_loc1053;
req  [19:0] cam_loc1054;
req  [19:0] cam_loc1055;
req  [19:0] cam_loc1056;
req  [19:0] cam_loc1057;
req  [19:0] cam_loc1058;
req  [19:0] cam_loc1059;
req  [19:0] cam_loc1060;
req  [19:0] cam_loc1061;
req  [19:0] cam_loc1062;
req  [19:0] cam_loc1063;
req  [19:0] cam_loc1064;
req  [19:0] cam_loc1065;
req  [19:0] cam_loc1066;
req  [19:0] cam_loc1067;
req  [19:0] cam_loc1068;
req  [19:0] cam_loc1069;
req  [19:0] cam_loc1070;
req  [19:0] cam_loc1071;
req  [19:0] cam_loc1072;
req  [19:0] cam_loc1073;
req  [19:0] cam_loc1074;
req  [19:0] cam_loc1075;
req  [19:0] cam_loc1076;
req  [19:0] cam_loc1077;
req  [19:0] cam_loc1078;
req  [19:0] cam_loc1079;
req  [19:0] cam_loc1080;
req  [19:0] cam_loc1081;
req  [19:0] cam_loc1082;
req  [19:0] cam_loc1083;
req  [19:0] cam_loc1084;
req  [19:0] cam_loc1085;
req  [19:0] cam_loc1086;
req  [19:0] cam_loc1087;
req  [19:0] cam_loc1088;
req  [19:0] cam_loc1089;
req  [19:0] cam_loc1090;
req  [19:0] cam_loc1091;
req  [19:0] cam_loc1092;
req  [19:0] cam_loc1093;
req  [19:0] cam_loc1094;
req  [19:0] cam_loc1095;
req  [19:0] cam_loc1096;
req  [19:0] cam_loc1097;
req  [19:0] cam_loc1098;
req  [19:0] cam_loc1099;

        always @ (posedge clk or negedge rst_an)
begin
if (!rst_an) begin
  wr_loc_counter <= 11+1'd0; // log2(CAMDEPTH) +1
       end else begin
  wr_loc_counter <= wr_location_counter[11] ? wr_location_counter : wr_location_counter + 1'b1;
       end
end
AH_srvfifo_11_CAMDEPTH u_wrloc_recirfifo (
.wr_valid(freeup_loc)
,.wr_ready(freedup_loc_valid)
,.wr_data(freedup_loc_ready)

,.rd_valid(recir_loc_valid)
,.rd_ready(recir_loc_ready)
,.rd_data(recir_loc)
);

assign internal_wr_en = wr_valid & (recir_loc_valid | ~wr_location_counter[11]);
assign internal_wr_ptr = ~wr_location_counter[11 + 1] ? ~wr_location_counter[10:0] : recir_loc;

assign wr_ready	= ~wr_location_counter[11 + 1] ? 1'b1 : recir_loc_valid;

assign recir_loc_ready	= ~wr_location_counter[11 + 1] ? 1'b0 : wr_valid;

always @ (posedge clk or negedge rst_an)
if (!rst_an) begin


	cam_loc0 <= 20'd0;
	cam_loc1 <= 20'd0;
	cam_loc2 <= 20'd0;
	cam_loc3 <= 20'd0;
	cam_loc4 <= 20'd0;
	cam_loc5 <= 20'd0;
	cam_loc6 <= 20'd0;
	cam_loc7 <= 20'd0;
	cam_loc8 <= 20'd0;
	cam_loc9 <= 20'd0;
	cam_loc10 <= 20'd0;
	cam_loc11 <= 20'd0;
	cam_loc12 <= 20'd0;
	cam_loc13 <= 20'd0;
	cam_loc14 <= 20'd0;
	cam_loc15 <= 20'd0;
	cam_loc16 <= 20'd0;
	cam_loc17 <= 20'd0;
	cam_loc18 <= 20'd0;
	cam_loc19 <= 20'd0;
	cam_loc20 <= 20'd0;
	cam_loc21 <= 20'd0;
	cam_loc22 <= 20'd0;
	cam_loc23 <= 20'd0;
	cam_loc24 <= 20'd0;
	cam_loc25 <= 20'd0;
	cam_loc26 <= 20'd0;
	cam_loc27 <= 20'd0;
	cam_loc28 <= 20'd0;
	cam_loc29 <= 20'd0;
	cam_loc30 <= 20'd0;
	cam_loc31 <= 20'd0;
	cam_loc32 <= 20'd0;
	cam_loc33 <= 20'd0;
	cam_loc34 <= 20'd0;
	cam_loc35 <= 20'd0;
	cam_loc36 <= 20'd0;
	cam_loc37 <= 20'd0;
	cam_loc38 <= 20'd0;
	cam_loc39 <= 20'd0;
	cam_loc40 <= 20'd0;
	cam_loc41 <= 20'd0;
	cam_loc42 <= 20'd0;
	cam_loc43 <= 20'd0;
	cam_loc44 <= 20'd0;
	cam_loc45 <= 20'd0;
	cam_loc46 <= 20'd0;
	cam_loc47 <= 20'd0;
	cam_loc48 <= 20'd0;
	cam_loc49 <= 20'd0;
	cam_loc50 <= 20'd0;
	cam_loc51 <= 20'd0;
	cam_loc52 <= 20'd0;
	cam_loc53 <= 20'd0;
	cam_loc54 <= 20'd0;
	cam_loc55 <= 20'd0;
	cam_loc56 <= 20'd0;
	cam_loc57 <= 20'd0;
	cam_loc58 <= 20'd0;
	cam_loc59 <= 20'd0;
	cam_loc60 <= 20'd0;
	cam_loc61 <= 20'd0;
	cam_loc62 <= 20'd0;
	cam_loc63 <= 20'd0;
	cam_loc64 <= 20'd0;
	cam_loc65 <= 20'd0;
	cam_loc66 <= 20'd0;
	cam_loc67 <= 20'd0;
	cam_loc68 <= 20'd0;
	cam_loc69 <= 20'd0;
	cam_loc70 <= 20'd0;
	cam_loc71 <= 20'd0;
	cam_loc72 <= 20'd0;
	cam_loc73 <= 20'd0;
	cam_loc74 <= 20'd0;
	cam_loc75 <= 20'd0;
	cam_loc76 <= 20'd0;
	cam_loc77 <= 20'd0;
	cam_loc78 <= 20'd0;
	cam_loc79 <= 20'd0;
	cam_loc80 <= 20'd0;
	cam_loc81 <= 20'd0;
	cam_loc82 <= 20'd0;
	cam_loc83 <= 20'd0;
	cam_loc84 <= 20'd0;
	cam_loc85 <= 20'd0;
	cam_loc86 <= 20'd0;
	cam_loc87 <= 20'd0;
	cam_loc88 <= 20'd0;
	cam_loc89 <= 20'd0;
	cam_loc90 <= 20'd0;
	cam_loc91 <= 20'd0;
	cam_loc92 <= 20'd0;
	cam_loc93 <= 20'd0;
	cam_loc94 <= 20'd0;
	cam_loc95 <= 20'd0;
	cam_loc96 <= 20'd0;
	cam_loc97 <= 20'd0;
	cam_loc98 <= 20'd0;
	cam_loc99 <= 20'd0;
	cam_loc100 <= 20'd0;
	cam_loc101 <= 20'd0;
	cam_loc102 <= 20'd0;
	cam_loc103 <= 20'd0;
	cam_loc104 <= 20'd0;
	cam_loc105 <= 20'd0;
	cam_loc106 <= 20'd0;
	cam_loc107 <= 20'd0;
	cam_loc108 <= 20'd0;
	cam_loc109 <= 20'd0;
	cam_loc110 <= 20'd0;
	cam_loc111 <= 20'd0;
	cam_loc112 <= 20'd0;
	cam_loc113 <= 20'd0;
	cam_loc114 <= 20'd0;
	cam_loc115 <= 20'd0;
	cam_loc116 <= 20'd0;
	cam_loc117 <= 20'd0;
	cam_loc118 <= 20'd0;
	cam_loc119 <= 20'd0;
	cam_loc120 <= 20'd0;
	cam_loc121 <= 20'd0;
	cam_loc122 <= 20'd0;
	cam_loc123 <= 20'd0;
	cam_loc124 <= 20'd0;
	cam_loc125 <= 20'd0;
	cam_loc126 <= 20'd0;
	cam_loc127 <= 20'd0;
	cam_loc128 <= 20'd0;
	cam_loc129 <= 20'd0;
	cam_loc130 <= 20'd0;
	cam_loc131 <= 20'd0;
	cam_loc132 <= 20'd0;
	cam_loc133 <= 20'd0;
	cam_loc134 <= 20'd0;
	cam_loc135 <= 20'd0;
	cam_loc136 <= 20'd0;
	cam_loc137 <= 20'd0;
	cam_loc138 <= 20'd0;
	cam_loc139 <= 20'd0;
	cam_loc140 <= 20'd0;
	cam_loc141 <= 20'd0;
	cam_loc142 <= 20'd0;
	cam_loc143 <= 20'd0;
	cam_loc144 <= 20'd0;
	cam_loc145 <= 20'd0;
	cam_loc146 <= 20'd0;
	cam_loc147 <= 20'd0;
	cam_loc148 <= 20'd0;
	cam_loc149 <= 20'd0;
	cam_loc150 <= 20'd0;
	cam_loc151 <= 20'd0;
	cam_loc152 <= 20'd0;
	cam_loc153 <= 20'd0;
	cam_loc154 <= 20'd0;
	cam_loc155 <= 20'd0;
	cam_loc156 <= 20'd0;
	cam_loc157 <= 20'd0;
	cam_loc158 <= 20'd0;
	cam_loc159 <= 20'd0;
	cam_loc160 <= 20'd0;
	cam_loc161 <= 20'd0;
	cam_loc162 <= 20'd0;
	cam_loc163 <= 20'd0;
	cam_loc164 <= 20'd0;
	cam_loc165 <= 20'd0;
	cam_loc166 <= 20'd0;
	cam_loc167 <= 20'd0;
	cam_loc168 <= 20'd0;
	cam_loc169 <= 20'd0;
	cam_loc170 <= 20'd0;
	cam_loc171 <= 20'd0;
	cam_loc172 <= 20'd0;
	cam_loc173 <= 20'd0;
	cam_loc174 <= 20'd0;
	cam_loc175 <= 20'd0;
	cam_loc176 <= 20'd0;
	cam_loc177 <= 20'd0;
	cam_loc178 <= 20'd0;
	cam_loc179 <= 20'd0;
	cam_loc180 <= 20'd0;
	cam_loc181 <= 20'd0;
	cam_loc182 <= 20'd0;
	cam_loc183 <= 20'd0;
	cam_loc184 <= 20'd0;
	cam_loc185 <= 20'd0;
	cam_loc186 <= 20'd0;
	cam_loc187 <= 20'd0;
	cam_loc188 <= 20'd0;
	cam_loc189 <= 20'd0;
	cam_loc190 <= 20'd0;
	cam_loc191 <= 20'd0;
	cam_loc192 <= 20'd0;
	cam_loc193 <= 20'd0;
	cam_loc194 <= 20'd0;
	cam_loc195 <= 20'd0;
	cam_loc196 <= 20'd0;
	cam_loc197 <= 20'd0;
	cam_loc198 <= 20'd0;
	cam_loc199 <= 20'd0;
	cam_loc200 <= 20'd0;
	cam_loc201 <= 20'd0;
	cam_loc202 <= 20'd0;
	cam_loc203 <= 20'd0;
	cam_loc204 <= 20'd0;
	cam_loc205 <= 20'd0;
	cam_loc206 <= 20'd0;
	cam_loc207 <= 20'd0;
	cam_loc208 <= 20'd0;
	cam_loc209 <= 20'd0;
	cam_loc210 <= 20'd0;
	cam_loc211 <= 20'd0;
	cam_loc212 <= 20'd0;
	cam_loc213 <= 20'd0;
	cam_loc214 <= 20'd0;
	cam_loc215 <= 20'd0;
	cam_loc216 <= 20'd0;
	cam_loc217 <= 20'd0;
	cam_loc218 <= 20'd0;
	cam_loc219 <= 20'd0;
	cam_loc220 <= 20'd0;
	cam_loc221 <= 20'd0;
	cam_loc222 <= 20'd0;
	cam_loc223 <= 20'd0;
	cam_loc224 <= 20'd0;
	cam_loc225 <= 20'd0;
	cam_loc226 <= 20'd0;
	cam_loc227 <= 20'd0;
	cam_loc228 <= 20'd0;
	cam_loc229 <= 20'd0;
	cam_loc230 <= 20'd0;
	cam_loc231 <= 20'd0;
	cam_loc232 <= 20'd0;
	cam_loc233 <= 20'd0;
	cam_loc234 <= 20'd0;
	cam_loc235 <= 20'd0;
	cam_loc236 <= 20'd0;
	cam_loc237 <= 20'd0;
	cam_loc238 <= 20'd0;
	cam_loc239 <= 20'd0;
	cam_loc240 <= 20'd0;
	cam_loc241 <= 20'd0;
	cam_loc242 <= 20'd0;
	cam_loc243 <= 20'd0;
	cam_loc244 <= 20'd0;
	cam_loc245 <= 20'd0;
	cam_loc246 <= 20'd0;
	cam_loc247 <= 20'd0;
	cam_loc248 <= 20'd0;
	cam_loc249 <= 20'd0;
	cam_loc250 <= 20'd0;
	cam_loc251 <= 20'd0;
	cam_loc252 <= 20'd0;
	cam_loc253 <= 20'd0;
	cam_loc254 <= 20'd0;
	cam_loc255 <= 20'd0;
	cam_loc256 <= 20'd0;
	cam_loc257 <= 20'd0;
	cam_loc258 <= 20'd0;
	cam_loc259 <= 20'd0;
	cam_loc260 <= 20'd0;
	cam_loc261 <= 20'd0;
	cam_loc262 <= 20'd0;
	cam_loc263 <= 20'd0;
	cam_loc264 <= 20'd0;
	cam_loc265 <= 20'd0;
	cam_loc266 <= 20'd0;
	cam_loc267 <= 20'd0;
	cam_loc268 <= 20'd0;
	cam_loc269 <= 20'd0;
	cam_loc270 <= 20'd0;
	cam_loc271 <= 20'd0;
	cam_loc272 <= 20'd0;
	cam_loc273 <= 20'd0;
	cam_loc274 <= 20'd0;
	cam_loc275 <= 20'd0;
	cam_loc276 <= 20'd0;
	cam_loc277 <= 20'd0;
	cam_loc278 <= 20'd0;
	cam_loc279 <= 20'd0;
	cam_loc280 <= 20'd0;
	cam_loc281 <= 20'd0;
	cam_loc282 <= 20'd0;
	cam_loc283 <= 20'd0;
	cam_loc284 <= 20'd0;
	cam_loc285 <= 20'd0;
	cam_loc286 <= 20'd0;
	cam_loc287 <= 20'd0;
	cam_loc288 <= 20'd0;
	cam_loc289 <= 20'd0;
	cam_loc290 <= 20'd0;
	cam_loc291 <= 20'd0;
	cam_loc292 <= 20'd0;
	cam_loc293 <= 20'd0;
	cam_loc294 <= 20'd0;
	cam_loc295 <= 20'd0;
	cam_loc296 <= 20'd0;
	cam_loc297 <= 20'd0;
	cam_loc298 <= 20'd0;
	cam_loc299 <= 20'd0;
	cam_loc300 <= 20'd0;
	cam_loc301 <= 20'd0;
	cam_loc302 <= 20'd0;
	cam_loc303 <= 20'd0;
	cam_loc304 <= 20'd0;
	cam_loc305 <= 20'd0;
	cam_loc306 <= 20'd0;
	cam_loc307 <= 20'd0;
	cam_loc308 <= 20'd0;
	cam_loc309 <= 20'd0;
	cam_loc310 <= 20'd0;
	cam_loc311 <= 20'd0;
	cam_loc312 <= 20'd0;
	cam_loc313 <= 20'd0;
	cam_loc314 <= 20'd0;
	cam_loc315 <= 20'd0;
	cam_loc316 <= 20'd0;
	cam_loc317 <= 20'd0;
	cam_loc318 <= 20'd0;
	cam_loc319 <= 20'd0;
	cam_loc320 <= 20'd0;
	cam_loc321 <= 20'd0;
	cam_loc322 <= 20'd0;
	cam_loc323 <= 20'd0;
	cam_loc324 <= 20'd0;
	cam_loc325 <= 20'd0;
	cam_loc326 <= 20'd0;
	cam_loc327 <= 20'd0;
	cam_loc328 <= 20'd0;
	cam_loc329 <= 20'd0;
	cam_loc330 <= 20'd0;
	cam_loc331 <= 20'd0;
	cam_loc332 <= 20'd0;
	cam_loc333 <= 20'd0;
	cam_loc334 <= 20'd0;
	cam_loc335 <= 20'd0;
	cam_loc336 <= 20'd0;
	cam_loc337 <= 20'd0;
	cam_loc338 <= 20'd0;
	cam_loc339 <= 20'd0;
	cam_loc340 <= 20'd0;
	cam_loc341 <= 20'd0;
	cam_loc342 <= 20'd0;
	cam_loc343 <= 20'd0;
	cam_loc344 <= 20'd0;
	cam_loc345 <= 20'd0;
	cam_loc346 <= 20'd0;
	cam_loc347 <= 20'd0;
	cam_loc348 <= 20'd0;
	cam_loc349 <= 20'd0;
	cam_loc350 <= 20'd0;
	cam_loc351 <= 20'd0;
	cam_loc352 <= 20'd0;
	cam_loc353 <= 20'd0;
	cam_loc354 <= 20'd0;
	cam_loc355 <= 20'd0;
	cam_loc356 <= 20'd0;
	cam_loc357 <= 20'd0;
	cam_loc358 <= 20'd0;
	cam_loc359 <= 20'd0;
	cam_loc360 <= 20'd0;
	cam_loc361 <= 20'd0;
	cam_loc362 <= 20'd0;
	cam_loc363 <= 20'd0;
	cam_loc364 <= 20'd0;
	cam_loc365 <= 20'd0;
	cam_loc366 <= 20'd0;
	cam_loc367 <= 20'd0;
	cam_loc368 <= 20'd0;
	cam_loc369 <= 20'd0;
	cam_loc370 <= 20'd0;
	cam_loc371 <= 20'd0;
	cam_loc372 <= 20'd0;
	cam_loc373 <= 20'd0;
	cam_loc374 <= 20'd0;
	cam_loc375 <= 20'd0;
	cam_loc376 <= 20'd0;
	cam_loc377 <= 20'd0;
	cam_loc378 <= 20'd0;
	cam_loc379 <= 20'd0;
	cam_loc380 <= 20'd0;
	cam_loc381 <= 20'd0;
	cam_loc382 <= 20'd0;
	cam_loc383 <= 20'd0;
	cam_loc384 <= 20'd0;
	cam_loc385 <= 20'd0;
	cam_loc386 <= 20'd0;
	cam_loc387 <= 20'd0;
	cam_loc388 <= 20'd0;
	cam_loc389 <= 20'd0;
	cam_loc390 <= 20'd0;
	cam_loc391 <= 20'd0;
	cam_loc392 <= 20'd0;
	cam_loc393 <= 20'd0;
	cam_loc394 <= 20'd0;
	cam_loc395 <= 20'd0;
	cam_loc396 <= 20'd0;
	cam_loc397 <= 20'd0;
	cam_loc398 <= 20'd0;
	cam_loc399 <= 20'd0;
	cam_loc400 <= 20'd0;
	cam_loc401 <= 20'd0;
	cam_loc402 <= 20'd0;
	cam_loc403 <= 20'd0;
	cam_loc404 <= 20'd0;
	cam_loc405 <= 20'd0;
	cam_loc406 <= 20'd0;
	cam_loc407 <= 20'd0;
	cam_loc408 <= 20'd0;
	cam_loc409 <= 20'd0;
	cam_loc410 <= 20'd0;
	cam_loc411 <= 20'd0;
	cam_loc412 <= 20'd0;
	cam_loc413 <= 20'd0;
	cam_loc414 <= 20'd0;
	cam_loc415 <= 20'd0;
	cam_loc416 <= 20'd0;
	cam_loc417 <= 20'd0;
	cam_loc418 <= 20'd0;
	cam_loc419 <= 20'd0;
	cam_loc420 <= 20'd0;
	cam_loc421 <= 20'd0;
	cam_loc422 <= 20'd0;
	cam_loc423 <= 20'd0;
	cam_loc424 <= 20'd0;
	cam_loc425 <= 20'd0;
	cam_loc426 <= 20'd0;
	cam_loc427 <= 20'd0;
	cam_loc428 <= 20'd0;
	cam_loc429 <= 20'd0;
	cam_loc430 <= 20'd0;
	cam_loc431 <= 20'd0;
	cam_loc432 <= 20'd0;
	cam_loc433 <= 20'd0;
	cam_loc434 <= 20'd0;
	cam_loc435 <= 20'd0;
	cam_loc436 <= 20'd0;
	cam_loc437 <= 20'd0;
	cam_loc438 <= 20'd0;
	cam_loc439 <= 20'd0;
	cam_loc440 <= 20'd0;
	cam_loc441 <= 20'd0;
	cam_loc442 <= 20'd0;
	cam_loc443 <= 20'd0;
	cam_loc444 <= 20'd0;
	cam_loc445 <= 20'd0;
	cam_loc446 <= 20'd0;
	cam_loc447 <= 20'd0;
	cam_loc448 <= 20'd0;
	cam_loc449 <= 20'd0;
	cam_loc450 <= 20'd0;
	cam_loc451 <= 20'd0;
	cam_loc452 <= 20'd0;
	cam_loc453 <= 20'd0;
	cam_loc454 <= 20'd0;
	cam_loc455 <= 20'd0;
	cam_loc456 <= 20'd0;
	cam_loc457 <= 20'd0;
	cam_loc458 <= 20'd0;
	cam_loc459 <= 20'd0;
	cam_loc460 <= 20'd0;
	cam_loc461 <= 20'd0;
	cam_loc462 <= 20'd0;
	cam_loc463 <= 20'd0;
	cam_loc464 <= 20'd0;
	cam_loc465 <= 20'd0;
	cam_loc466 <= 20'd0;
	cam_loc467 <= 20'd0;
	cam_loc468 <= 20'd0;
	cam_loc469 <= 20'd0;
	cam_loc470 <= 20'd0;
	cam_loc471 <= 20'd0;
	cam_loc472 <= 20'd0;
	cam_loc473 <= 20'd0;
	cam_loc474 <= 20'd0;
	cam_loc475 <= 20'd0;
	cam_loc476 <= 20'd0;
	cam_loc477 <= 20'd0;
	cam_loc478 <= 20'd0;
	cam_loc479 <= 20'd0;
	cam_loc480 <= 20'd0;
	cam_loc481 <= 20'd0;
	cam_loc482 <= 20'd0;
	cam_loc483 <= 20'd0;
	cam_loc484 <= 20'd0;
	cam_loc485 <= 20'd0;
	cam_loc486 <= 20'd0;
	cam_loc487 <= 20'd0;
	cam_loc488 <= 20'd0;
	cam_loc489 <= 20'd0;
	cam_loc490 <= 20'd0;
	cam_loc491 <= 20'd0;
	cam_loc492 <= 20'd0;
	cam_loc493 <= 20'd0;
	cam_loc494 <= 20'd0;
	cam_loc495 <= 20'd0;
	cam_loc496 <= 20'd0;
	cam_loc497 <= 20'd0;
	cam_loc498 <= 20'd0;
	cam_loc499 <= 20'd0;
	cam_loc500 <= 20'd0;
	cam_loc501 <= 20'd0;
	cam_loc502 <= 20'd0;
	cam_loc503 <= 20'd0;
	cam_loc504 <= 20'd0;
	cam_loc505 <= 20'd0;
	cam_loc506 <= 20'd0;
	cam_loc507 <= 20'd0;
	cam_loc508 <= 20'd0;
	cam_loc509 <= 20'd0;
	cam_loc510 <= 20'd0;
	cam_loc511 <= 20'd0;
	cam_loc512 <= 20'd0;
	cam_loc513 <= 20'd0;
	cam_loc514 <= 20'd0;
	cam_loc515 <= 20'd0;
	cam_loc516 <= 20'd0;
	cam_loc517 <= 20'd0;
	cam_loc518 <= 20'd0;
	cam_loc519 <= 20'd0;
	cam_loc520 <= 20'd0;
	cam_loc521 <= 20'd0;
	cam_loc522 <= 20'd0;
	cam_loc523 <= 20'd0;
	cam_loc524 <= 20'd0;
	cam_loc525 <= 20'd0;
	cam_loc526 <= 20'd0;
	cam_loc527 <= 20'd0;
	cam_loc528 <= 20'd0;
	cam_loc529 <= 20'd0;
	cam_loc530 <= 20'd0;
	cam_loc531 <= 20'd0;
	cam_loc532 <= 20'd0;
	cam_loc533 <= 20'd0;
	cam_loc534 <= 20'd0;
	cam_loc535 <= 20'd0;
	cam_loc536 <= 20'd0;
	cam_loc537 <= 20'd0;
	cam_loc538 <= 20'd0;
	cam_loc539 <= 20'd0;
	cam_loc540 <= 20'd0;
	cam_loc541 <= 20'd0;
	cam_loc542 <= 20'd0;
	cam_loc543 <= 20'd0;
	cam_loc544 <= 20'd0;
	cam_loc545 <= 20'd0;
	cam_loc546 <= 20'd0;
	cam_loc547 <= 20'd0;
	cam_loc548 <= 20'd0;
	cam_loc549 <= 20'd0;
	cam_loc550 <= 20'd0;
	cam_loc551 <= 20'd0;
	cam_loc552 <= 20'd0;
	cam_loc553 <= 20'd0;
	cam_loc554 <= 20'd0;
	cam_loc555 <= 20'd0;
	cam_loc556 <= 20'd0;
	cam_loc557 <= 20'd0;
	cam_loc558 <= 20'd0;
	cam_loc559 <= 20'd0;
	cam_loc560 <= 20'd0;
	cam_loc561 <= 20'd0;
	cam_loc562 <= 20'd0;
	cam_loc563 <= 20'd0;
	cam_loc564 <= 20'd0;
	cam_loc565 <= 20'd0;
	cam_loc566 <= 20'd0;
	cam_loc567 <= 20'd0;
	cam_loc568 <= 20'd0;
	cam_loc569 <= 20'd0;
	cam_loc570 <= 20'd0;
	cam_loc571 <= 20'd0;
	cam_loc572 <= 20'd0;
	cam_loc573 <= 20'd0;
	cam_loc574 <= 20'd0;
	cam_loc575 <= 20'd0;
	cam_loc576 <= 20'd0;
	cam_loc577 <= 20'd0;
	cam_loc578 <= 20'd0;
	cam_loc579 <= 20'd0;
	cam_loc580 <= 20'd0;
	cam_loc581 <= 20'd0;
	cam_loc582 <= 20'd0;
	cam_loc583 <= 20'd0;
	cam_loc584 <= 20'd0;
	cam_loc585 <= 20'd0;
	cam_loc586 <= 20'd0;
	cam_loc587 <= 20'd0;
	cam_loc588 <= 20'd0;
	cam_loc589 <= 20'd0;
	cam_loc590 <= 20'd0;
	cam_loc591 <= 20'd0;
	cam_loc592 <= 20'd0;
	cam_loc593 <= 20'd0;
	cam_loc594 <= 20'd0;
	cam_loc595 <= 20'd0;
	cam_loc596 <= 20'd0;
	cam_loc597 <= 20'd0;
	cam_loc598 <= 20'd0;
	cam_loc599 <= 20'd0;
	cam_loc600 <= 20'd0;
	cam_loc601 <= 20'd0;
	cam_loc602 <= 20'd0;
	cam_loc603 <= 20'd0;
	cam_loc604 <= 20'd0;
	cam_loc605 <= 20'd0;
	cam_loc606 <= 20'd0;
	cam_loc607 <= 20'd0;
	cam_loc608 <= 20'd0;
	cam_loc609 <= 20'd0;
	cam_loc610 <= 20'd0;
	cam_loc611 <= 20'd0;
	cam_loc612 <= 20'd0;
	cam_loc613 <= 20'd0;
	cam_loc614 <= 20'd0;
	cam_loc615 <= 20'd0;
	cam_loc616 <= 20'd0;
	cam_loc617 <= 20'd0;
	cam_loc618 <= 20'd0;
	cam_loc619 <= 20'd0;
	cam_loc620 <= 20'd0;
	cam_loc621 <= 20'd0;
	cam_loc622 <= 20'd0;
	cam_loc623 <= 20'd0;
	cam_loc624 <= 20'd0;
	cam_loc625 <= 20'd0;
	cam_loc626 <= 20'd0;
	cam_loc627 <= 20'd0;
	cam_loc628 <= 20'd0;
	cam_loc629 <= 20'd0;
	cam_loc630 <= 20'd0;
	cam_loc631 <= 20'd0;
	cam_loc632 <= 20'd0;
	cam_loc633 <= 20'd0;
	cam_loc634 <= 20'd0;
	cam_loc635 <= 20'd0;
	cam_loc636 <= 20'd0;
	cam_loc637 <= 20'd0;
	cam_loc638 <= 20'd0;
	cam_loc639 <= 20'd0;
	cam_loc640 <= 20'd0;
	cam_loc641 <= 20'd0;
	cam_loc642 <= 20'd0;
	cam_loc643 <= 20'd0;
	cam_loc644 <= 20'd0;
	cam_loc645 <= 20'd0;
	cam_loc646 <= 20'd0;
	cam_loc647 <= 20'd0;
	cam_loc648 <= 20'd0;
	cam_loc649 <= 20'd0;
	cam_loc650 <= 20'd0;
	cam_loc651 <= 20'd0;
	cam_loc652 <= 20'd0;
	cam_loc653 <= 20'd0;
	cam_loc654 <= 20'd0;
	cam_loc655 <= 20'd0;
	cam_loc656 <= 20'd0;
	cam_loc657 <= 20'd0;
	cam_loc658 <= 20'd0;
	cam_loc659 <= 20'd0;
	cam_loc660 <= 20'd0;
	cam_loc661 <= 20'd0;
	cam_loc662 <= 20'd0;
	cam_loc663 <= 20'd0;
	cam_loc664 <= 20'd0;
	cam_loc665 <= 20'd0;
	cam_loc666 <= 20'd0;
	cam_loc667 <= 20'd0;
	cam_loc668 <= 20'd0;
	cam_loc669 <= 20'd0;
	cam_loc670 <= 20'd0;
	cam_loc671 <= 20'd0;
	cam_loc672 <= 20'd0;
	cam_loc673 <= 20'd0;
	cam_loc674 <= 20'd0;
	cam_loc675 <= 20'd0;
	cam_loc676 <= 20'd0;
	cam_loc677 <= 20'd0;
	cam_loc678 <= 20'd0;
	cam_loc679 <= 20'd0;
	cam_loc680 <= 20'd0;
	cam_loc681 <= 20'd0;
	cam_loc682 <= 20'd0;
	cam_loc683 <= 20'd0;
	cam_loc684 <= 20'd0;
	cam_loc685 <= 20'd0;
	cam_loc686 <= 20'd0;
	cam_loc687 <= 20'd0;
	cam_loc688 <= 20'd0;
	cam_loc689 <= 20'd0;
	cam_loc690 <= 20'd0;
	cam_loc691 <= 20'd0;
	cam_loc692 <= 20'd0;
	cam_loc693 <= 20'd0;
	cam_loc694 <= 20'd0;
	cam_loc695 <= 20'd0;
	cam_loc696 <= 20'd0;
	cam_loc697 <= 20'd0;
	cam_loc698 <= 20'd0;
	cam_loc699 <= 20'd0;
	cam_loc700 <= 20'd0;
	cam_loc701 <= 20'd0;
	cam_loc702 <= 20'd0;
	cam_loc703 <= 20'd0;
	cam_loc704 <= 20'd0;
	cam_loc705 <= 20'd0;
	cam_loc706 <= 20'd0;
	cam_loc707 <= 20'd0;
	cam_loc708 <= 20'd0;
	cam_loc709 <= 20'd0;
	cam_loc710 <= 20'd0;
	cam_loc711 <= 20'd0;
	cam_loc712 <= 20'd0;
	cam_loc713 <= 20'd0;
	cam_loc714 <= 20'd0;
	cam_loc715 <= 20'd0;
	cam_loc716 <= 20'd0;
	cam_loc717 <= 20'd0;
	cam_loc718 <= 20'd0;
	cam_loc719 <= 20'd0;
	cam_loc720 <= 20'd0;
	cam_loc721 <= 20'd0;
	cam_loc722 <= 20'd0;
	cam_loc723 <= 20'd0;
	cam_loc724 <= 20'd0;
	cam_loc725 <= 20'd0;
	cam_loc726 <= 20'd0;
	cam_loc727 <= 20'd0;
	cam_loc728 <= 20'd0;
	cam_loc729 <= 20'd0;
	cam_loc730 <= 20'd0;
	cam_loc731 <= 20'd0;
	cam_loc732 <= 20'd0;
	cam_loc733 <= 20'd0;
	cam_loc734 <= 20'd0;
	cam_loc735 <= 20'd0;
	cam_loc736 <= 20'd0;
	cam_loc737 <= 20'd0;
	cam_loc738 <= 20'd0;
	cam_loc739 <= 20'd0;
	cam_loc740 <= 20'd0;
	cam_loc741 <= 20'd0;
	cam_loc742 <= 20'd0;
	cam_loc743 <= 20'd0;
	cam_loc744 <= 20'd0;
	cam_loc745 <= 20'd0;
	cam_loc746 <= 20'd0;
	cam_loc747 <= 20'd0;
	cam_loc748 <= 20'd0;
	cam_loc749 <= 20'd0;
	cam_loc750 <= 20'd0;
	cam_loc751 <= 20'd0;
	cam_loc752 <= 20'd0;
	cam_loc753 <= 20'd0;
	cam_loc754 <= 20'd0;
	cam_loc755 <= 20'd0;
	cam_loc756 <= 20'd0;
	cam_loc757 <= 20'd0;
	cam_loc758 <= 20'd0;
	cam_loc759 <= 20'd0;
	cam_loc760 <= 20'd0;
	cam_loc761 <= 20'd0;
	cam_loc762 <= 20'd0;
	cam_loc763 <= 20'd0;
	cam_loc764 <= 20'd0;
	cam_loc765 <= 20'd0;
	cam_loc766 <= 20'd0;
	cam_loc767 <= 20'd0;
	cam_loc768 <= 20'd0;
	cam_loc769 <= 20'd0;
	cam_loc770 <= 20'd0;
	cam_loc771 <= 20'd0;
	cam_loc772 <= 20'd0;
	cam_loc773 <= 20'd0;
	cam_loc774 <= 20'd0;
	cam_loc775 <= 20'd0;
	cam_loc776 <= 20'd0;
	cam_loc777 <= 20'd0;
	cam_loc778 <= 20'd0;
	cam_loc779 <= 20'd0;
	cam_loc780 <= 20'd0;
	cam_loc781 <= 20'd0;
	cam_loc782 <= 20'd0;
	cam_loc783 <= 20'd0;
	cam_loc784 <= 20'd0;
	cam_loc785 <= 20'd0;
	cam_loc786 <= 20'd0;
	cam_loc787 <= 20'd0;
	cam_loc788 <= 20'd0;
	cam_loc789 <= 20'd0;
	cam_loc790 <= 20'd0;
	cam_loc791 <= 20'd0;
	cam_loc792 <= 20'd0;
	cam_loc793 <= 20'd0;
	cam_loc794 <= 20'd0;
	cam_loc795 <= 20'd0;
	cam_loc796 <= 20'd0;
	cam_loc797 <= 20'd0;
	cam_loc798 <= 20'd0;
	cam_loc799 <= 20'd0;
	cam_loc800 <= 20'd0;
	cam_loc801 <= 20'd0;
	cam_loc802 <= 20'd0;
	cam_loc803 <= 20'd0;
	cam_loc804 <= 20'd0;
	cam_loc805 <= 20'd0;
	cam_loc806 <= 20'd0;
	cam_loc807 <= 20'd0;
	cam_loc808 <= 20'd0;
	cam_loc809 <= 20'd0;
	cam_loc810 <= 20'd0;
	cam_loc811 <= 20'd0;
	cam_loc812 <= 20'd0;
	cam_loc813 <= 20'd0;
	cam_loc814 <= 20'd0;
	cam_loc815 <= 20'd0;
	cam_loc816 <= 20'd0;
	cam_loc817 <= 20'd0;
	cam_loc818 <= 20'd0;
	cam_loc819 <= 20'd0;
	cam_loc820 <= 20'd0;
	cam_loc821 <= 20'd0;
	cam_loc822 <= 20'd0;
	cam_loc823 <= 20'd0;
	cam_loc824 <= 20'd0;
	cam_loc825 <= 20'd0;
	cam_loc826 <= 20'd0;
	cam_loc827 <= 20'd0;
	cam_loc828 <= 20'd0;
	cam_loc829 <= 20'd0;
	cam_loc830 <= 20'd0;
	cam_loc831 <= 20'd0;
	cam_loc832 <= 20'd0;
	cam_loc833 <= 20'd0;
	cam_loc834 <= 20'd0;
	cam_loc835 <= 20'd0;
	cam_loc836 <= 20'd0;
	cam_loc837 <= 20'd0;
	cam_loc838 <= 20'd0;
	cam_loc839 <= 20'd0;
	cam_loc840 <= 20'd0;
	cam_loc841 <= 20'd0;
	cam_loc842 <= 20'd0;
	cam_loc843 <= 20'd0;
	cam_loc844 <= 20'd0;
	cam_loc845 <= 20'd0;
	cam_loc846 <= 20'd0;
	cam_loc847 <= 20'd0;
	cam_loc848 <= 20'd0;
	cam_loc849 <= 20'd0;
	cam_loc850 <= 20'd0;
	cam_loc851 <= 20'd0;
	cam_loc852 <= 20'd0;
	cam_loc853 <= 20'd0;
	cam_loc854 <= 20'd0;
	cam_loc855 <= 20'd0;
	cam_loc856 <= 20'd0;
	cam_loc857 <= 20'd0;
	cam_loc858 <= 20'd0;
	cam_loc859 <= 20'd0;
	cam_loc860 <= 20'd0;
	cam_loc861 <= 20'd0;
	cam_loc862 <= 20'd0;
	cam_loc863 <= 20'd0;
	cam_loc864 <= 20'd0;
	cam_loc865 <= 20'd0;
	cam_loc866 <= 20'd0;
	cam_loc867 <= 20'd0;
	cam_loc868 <= 20'd0;
	cam_loc869 <= 20'd0;
	cam_loc870 <= 20'd0;
	cam_loc871 <= 20'd0;
	cam_loc872 <= 20'd0;
	cam_loc873 <= 20'd0;
	cam_loc874 <= 20'd0;
	cam_loc875 <= 20'd0;
	cam_loc876 <= 20'd0;
	cam_loc877 <= 20'd0;
	cam_loc878 <= 20'd0;
	cam_loc879 <= 20'd0;
	cam_loc880 <= 20'd0;
	cam_loc881 <= 20'd0;
	cam_loc882 <= 20'd0;
	cam_loc883 <= 20'd0;
	cam_loc884 <= 20'd0;
	cam_loc885 <= 20'd0;
	cam_loc886 <= 20'd0;
	cam_loc887 <= 20'd0;
	cam_loc888 <= 20'd0;
	cam_loc889 <= 20'd0;
	cam_loc890 <= 20'd0;
	cam_loc891 <= 20'd0;
	cam_loc892 <= 20'd0;
	cam_loc893 <= 20'd0;
	cam_loc894 <= 20'd0;
	cam_loc895 <= 20'd0;
	cam_loc896 <= 20'd0;
	cam_loc897 <= 20'd0;
	cam_loc898 <= 20'd0;
	cam_loc899 <= 20'd0;
	cam_loc900 <= 20'd0;
	cam_loc901 <= 20'd0;
	cam_loc902 <= 20'd0;
	cam_loc903 <= 20'd0;
	cam_loc904 <= 20'd0;
	cam_loc905 <= 20'd0;
	cam_loc906 <= 20'd0;
	cam_loc907 <= 20'd0;
	cam_loc908 <= 20'd0;
	cam_loc909 <= 20'd0;
	cam_loc910 <= 20'd0;
	cam_loc911 <= 20'd0;
	cam_loc912 <= 20'd0;
	cam_loc913 <= 20'd0;
	cam_loc914 <= 20'd0;
	cam_loc915 <= 20'd0;
	cam_loc916 <= 20'd0;
	cam_loc917 <= 20'd0;
	cam_loc918 <= 20'd0;
	cam_loc919 <= 20'd0;
	cam_loc920 <= 20'd0;
	cam_loc921 <= 20'd0;
	cam_loc922 <= 20'd0;
	cam_loc923 <= 20'd0;
	cam_loc924 <= 20'd0;
	cam_loc925 <= 20'd0;
	cam_loc926 <= 20'd0;
	cam_loc927 <= 20'd0;
	cam_loc928 <= 20'd0;
	cam_loc929 <= 20'd0;
	cam_loc930 <= 20'd0;
	cam_loc931 <= 20'd0;
	cam_loc932 <= 20'd0;
	cam_loc933 <= 20'd0;
	cam_loc934 <= 20'd0;
	cam_loc935 <= 20'd0;
	cam_loc936 <= 20'd0;
	cam_loc937 <= 20'd0;
	cam_loc938 <= 20'd0;
	cam_loc939 <= 20'd0;
	cam_loc940 <= 20'd0;
	cam_loc941 <= 20'd0;
	cam_loc942 <= 20'd0;
	cam_loc943 <= 20'd0;
	cam_loc944 <= 20'd0;
	cam_loc945 <= 20'd0;
	cam_loc946 <= 20'd0;
	cam_loc947 <= 20'd0;
	cam_loc948 <= 20'd0;
	cam_loc949 <= 20'd0;
	cam_loc950 <= 20'd0;
	cam_loc951 <= 20'd0;
	cam_loc952 <= 20'd0;
	cam_loc953 <= 20'd0;
	cam_loc954 <= 20'd0;
	cam_loc955 <= 20'd0;
	cam_loc956 <= 20'd0;
	cam_loc957 <= 20'd0;
	cam_loc958 <= 20'd0;
	cam_loc959 <= 20'd0;
	cam_loc960 <= 20'd0;
	cam_loc961 <= 20'd0;
	cam_loc962 <= 20'd0;
	cam_loc963 <= 20'd0;
	cam_loc964 <= 20'd0;
	cam_loc965 <= 20'd0;
	cam_loc966 <= 20'd0;
	cam_loc967 <= 20'd0;
	cam_loc968 <= 20'd0;
	cam_loc969 <= 20'd0;
	cam_loc970 <= 20'd0;
	cam_loc971 <= 20'd0;
	cam_loc972 <= 20'd0;
	cam_loc973 <= 20'd0;
	cam_loc974 <= 20'd0;
	cam_loc975 <= 20'd0;
	cam_loc976 <= 20'd0;
	cam_loc977 <= 20'd0;
	cam_loc978 <= 20'd0;
	cam_loc979 <= 20'd0;
	cam_loc980 <= 20'd0;
	cam_loc981 <= 20'd0;
	cam_loc982 <= 20'd0;
	cam_loc983 <= 20'd0;
	cam_loc984 <= 20'd0;
	cam_loc985 <= 20'd0;
	cam_loc986 <= 20'd0;
	cam_loc987 <= 20'd0;
	cam_loc988 <= 20'd0;
	cam_loc989 <= 20'd0;
	cam_loc990 <= 20'd0;
	cam_loc991 <= 20'd0;
	cam_loc992 <= 20'd0;
	cam_loc993 <= 20'd0;
	cam_loc994 <= 20'd0;
	cam_loc995 <= 20'd0;
	cam_loc996 <= 20'd0;
	cam_loc997 <= 20'd0;
	cam_loc998 <= 20'd0;
	cam_loc999 <= 20'd0;
	cam_loc1000 <= 20'd0;
	cam_loc1001 <= 20'd0;
	cam_loc1002 <= 20'd0;
	cam_loc1003 <= 20'd0;
	cam_loc1004 <= 20'd0;
	cam_loc1005 <= 20'd0;
	cam_loc1006 <= 20'd0;
	cam_loc1007 <= 20'd0;
	cam_loc1008 <= 20'd0;
	cam_loc1009 <= 20'd0;
	cam_loc1010 <= 20'd0;
	cam_loc1011 <= 20'd0;
	cam_loc1012 <= 20'd0;
	cam_loc1013 <= 20'd0;
	cam_loc1014 <= 20'd0;
	cam_loc1015 <= 20'd0;
	cam_loc1016 <= 20'd0;
	cam_loc1017 <= 20'd0;
	cam_loc1018 <= 20'd0;
	cam_loc1019 <= 20'd0;
	cam_loc1020 <= 20'd0;
	cam_loc1021 <= 20'd0;
	cam_loc1022 <= 20'd0;
	cam_loc1023 <= 20'd0;
	cam_loc1024 <= 20'd0;
	cam_loc1025 <= 20'd0;
	cam_loc1026 <= 20'd0;
	cam_loc1027 <= 20'd0;
	cam_loc1028 <= 20'd0;
	cam_loc1029 <= 20'd0;
	cam_loc1030 <= 20'd0;
	cam_loc1031 <= 20'd0;
	cam_loc1032 <= 20'd0;
	cam_loc1033 <= 20'd0;
	cam_loc1034 <= 20'd0;
	cam_loc1035 <= 20'd0;
	cam_loc1036 <= 20'd0;
	cam_loc1037 <= 20'd0;
	cam_loc1038 <= 20'd0;
	cam_loc1039 <= 20'd0;
	cam_loc1040 <= 20'd0;
	cam_loc1041 <= 20'd0;
	cam_loc1042 <= 20'd0;
	cam_loc1043 <= 20'd0;
	cam_loc1044 <= 20'd0;
	cam_loc1045 <= 20'd0;
	cam_loc1046 <= 20'd0;
	cam_loc1047 <= 20'd0;
	cam_loc1048 <= 20'd0;
	cam_loc1049 <= 20'd0;
	cam_loc1050 <= 20'd0;
	cam_loc1051 <= 20'd0;
	cam_loc1052 <= 20'd0;
	cam_loc1053 <= 20'd0;
	cam_loc1054 <= 20'd0;
	cam_loc1055 <= 20'd0;
	cam_loc1056 <= 20'd0;
	cam_loc1057 <= 20'd0;
	cam_loc1058 <= 20'd0;
	cam_loc1059 <= 20'd0;
	cam_loc1060 <= 20'd0;
	cam_loc1061 <= 20'd0;
	cam_loc1062 <= 20'd0;
	cam_loc1063 <= 20'd0;
	cam_loc1064 <= 20'd0;
	cam_loc1065 <= 20'd0;
	cam_loc1066 <= 20'd0;
	cam_loc1067 <= 20'd0;
	cam_loc1068 <= 20'd0;
	cam_loc1069 <= 20'd0;
	cam_loc1070 <= 20'd0;
	cam_loc1071 <= 20'd0;
	cam_loc1072 <= 20'd0;
	cam_loc1073 <= 20'd0;
	cam_loc1074 <= 20'd0;
	cam_loc1075 <= 20'd0;
	cam_loc1076 <= 20'd0;
	cam_loc1077 <= 20'd0;
	cam_loc1078 <= 20'd0;
	cam_loc1079 <= 20'd0;
	cam_loc1080 <= 20'd0;
	cam_loc1081 <= 20'd0;
	cam_loc1082 <= 20'd0;
	cam_loc1083 <= 20'd0;
	cam_loc1084 <= 20'd0;
	cam_loc1085 <= 20'd0;
	cam_loc1086 <= 20'd0;
	cam_loc1087 <= 20'd0;
	cam_loc1088 <= 20'd0;
	cam_loc1089 <= 20'd0;
	cam_loc1090 <= 20'd0;
	cam_loc1091 <= 20'd0;
	cam_loc1092 <= 20'd0;
	cam_loc1093 <= 20'd0;
	cam_loc1094 <= 20'd0;
	cam_loc1095 <= 20'd0;
	cam_loc1096 <= 20'd0;
	cam_loc1097 <= 20'd0;
	cam_loc1098 <= 20'd0;
	cam_loc1099 <= 20'd0;


end else begin

	cam_loc0 <= (internal_wr_en & (internal_wr_ptr == 11'd0) ) ? wr_data : cam_loc0;
	cam_loc1 <= (internal_wr_en & (internal_wr_ptr == 11'd1) ) ? wr_data : cam_loc1;
	cam_loc2 <= (internal_wr_en & (internal_wr_ptr == 11'd2) ) ? wr_data : cam_loc2;
	cam_loc3 <= (internal_wr_en & (internal_wr_ptr == 11'd3) ) ? wr_data : cam_loc3;
	cam_loc4 <= (internal_wr_en & (internal_wr_ptr == 11'd4) ) ? wr_data : cam_loc4;
	cam_loc5 <= (internal_wr_en & (internal_wr_ptr == 11'd5) ) ? wr_data : cam_loc5;
	cam_loc6 <= (internal_wr_en & (internal_wr_ptr == 11'd6) ) ? wr_data : cam_loc6;
	cam_loc7 <= (internal_wr_en & (internal_wr_ptr == 11'd7) ) ? wr_data : cam_loc7;
	cam_loc8 <= (internal_wr_en & (internal_wr_ptr == 11'd8) ) ? wr_data : cam_loc8;
	cam_loc9 <= (internal_wr_en & (internal_wr_ptr == 11'd9) ) ? wr_data : cam_loc9;
	cam_loc10 <= (internal_wr_en & (internal_wr_ptr == 11'd10) ) ? wr_data : cam_loc10;
	cam_loc11 <= (internal_wr_en & (internal_wr_ptr == 11'd11) ) ? wr_data : cam_loc11;
	cam_loc12 <= (internal_wr_en & (internal_wr_ptr == 11'd12) ) ? wr_data : cam_loc12;
	cam_loc13 <= (internal_wr_en & (internal_wr_ptr == 11'd13) ) ? wr_data : cam_loc13;
	cam_loc14 <= (internal_wr_en & (internal_wr_ptr == 11'd14) ) ? wr_data : cam_loc14;
	cam_loc15 <= (internal_wr_en & (internal_wr_ptr == 11'd15) ) ? wr_data : cam_loc15;
	cam_loc16 <= (internal_wr_en & (internal_wr_ptr == 11'd16) ) ? wr_data : cam_loc16;
	cam_loc17 <= (internal_wr_en & (internal_wr_ptr == 11'd17) ) ? wr_data : cam_loc17;
	cam_loc18 <= (internal_wr_en & (internal_wr_ptr == 11'd18) ) ? wr_data : cam_loc18;
	cam_loc19 <= (internal_wr_en & (internal_wr_ptr == 11'd19) ) ? wr_data : cam_loc19;
	cam_loc20 <= (internal_wr_en & (internal_wr_ptr == 11'd20) ) ? wr_data : cam_loc20;
	cam_loc21 <= (internal_wr_en & (internal_wr_ptr == 11'd21) ) ? wr_data : cam_loc21;
	cam_loc22 <= (internal_wr_en & (internal_wr_ptr == 11'd22) ) ? wr_data : cam_loc22;
	cam_loc23 <= (internal_wr_en & (internal_wr_ptr == 11'd23) ) ? wr_data : cam_loc23;
	cam_loc24 <= (internal_wr_en & (internal_wr_ptr == 11'd24) ) ? wr_data : cam_loc24;
	cam_loc25 <= (internal_wr_en & (internal_wr_ptr == 11'd25) ) ? wr_data : cam_loc25;
	cam_loc26 <= (internal_wr_en & (internal_wr_ptr == 11'd26) ) ? wr_data : cam_loc26;
	cam_loc27 <= (internal_wr_en & (internal_wr_ptr == 11'd27) ) ? wr_data : cam_loc27;
	cam_loc28 <= (internal_wr_en & (internal_wr_ptr == 11'd28) ) ? wr_data : cam_loc28;
	cam_loc29 <= (internal_wr_en & (internal_wr_ptr == 11'd29) ) ? wr_data : cam_loc29;
	cam_loc30 <= (internal_wr_en & (internal_wr_ptr == 11'd30) ) ? wr_data : cam_loc30;
	cam_loc31 <= (internal_wr_en & (internal_wr_ptr == 11'd31) ) ? wr_data : cam_loc31;
	cam_loc32 <= (internal_wr_en & (internal_wr_ptr == 11'd32) ) ? wr_data : cam_loc32;
	cam_loc33 <= (internal_wr_en & (internal_wr_ptr == 11'd33) ) ? wr_data : cam_loc33;
	cam_loc34 <= (internal_wr_en & (internal_wr_ptr == 11'd34) ) ? wr_data : cam_loc34;
	cam_loc35 <= (internal_wr_en & (internal_wr_ptr == 11'd35) ) ? wr_data : cam_loc35;
	cam_loc36 <= (internal_wr_en & (internal_wr_ptr == 11'd36) ) ? wr_data : cam_loc36;
	cam_loc37 <= (internal_wr_en & (internal_wr_ptr == 11'd37) ) ? wr_data : cam_loc37;
	cam_loc38 <= (internal_wr_en & (internal_wr_ptr == 11'd38) ) ? wr_data : cam_loc38;
	cam_loc39 <= (internal_wr_en & (internal_wr_ptr == 11'd39) ) ? wr_data : cam_loc39;
	cam_loc40 <= (internal_wr_en & (internal_wr_ptr == 11'd40) ) ? wr_data : cam_loc40;
	cam_loc41 <= (internal_wr_en & (internal_wr_ptr == 11'd41) ) ? wr_data : cam_loc41;
	cam_loc42 <= (internal_wr_en & (internal_wr_ptr == 11'd42) ) ? wr_data : cam_loc42;
	cam_loc43 <= (internal_wr_en & (internal_wr_ptr == 11'd43) ) ? wr_data : cam_loc43;
	cam_loc44 <= (internal_wr_en & (internal_wr_ptr == 11'd44) ) ? wr_data : cam_loc44;
	cam_loc45 <= (internal_wr_en & (internal_wr_ptr == 11'd45) ) ? wr_data : cam_loc45;
	cam_loc46 <= (internal_wr_en & (internal_wr_ptr == 11'd46) ) ? wr_data : cam_loc46;
	cam_loc47 <= (internal_wr_en & (internal_wr_ptr == 11'd47) ) ? wr_data : cam_loc47;
	cam_loc48 <= (internal_wr_en & (internal_wr_ptr == 11'd48) ) ? wr_data : cam_loc48;
	cam_loc49 <= (internal_wr_en & (internal_wr_ptr == 11'd49) ) ? wr_data : cam_loc49;
	cam_loc50 <= (internal_wr_en & (internal_wr_ptr == 11'd50) ) ? wr_data : cam_loc50;
	cam_loc51 <= (internal_wr_en & (internal_wr_ptr == 11'd51) ) ? wr_data : cam_loc51;
	cam_loc52 <= (internal_wr_en & (internal_wr_ptr == 11'd52) ) ? wr_data : cam_loc52;
	cam_loc53 <= (internal_wr_en & (internal_wr_ptr == 11'd53) ) ? wr_data : cam_loc53;
	cam_loc54 <= (internal_wr_en & (internal_wr_ptr == 11'd54) ) ? wr_data : cam_loc54;
	cam_loc55 <= (internal_wr_en & (internal_wr_ptr == 11'd55) ) ? wr_data : cam_loc55;
	cam_loc56 <= (internal_wr_en & (internal_wr_ptr == 11'd56) ) ? wr_data : cam_loc56;
	cam_loc57 <= (internal_wr_en & (internal_wr_ptr == 11'd57) ) ? wr_data : cam_loc57;
	cam_loc58 <= (internal_wr_en & (internal_wr_ptr == 11'd58) ) ? wr_data : cam_loc58;
	cam_loc59 <= (internal_wr_en & (internal_wr_ptr == 11'd59) ) ? wr_data : cam_loc59;
	cam_loc60 <= (internal_wr_en & (internal_wr_ptr == 11'd60) ) ? wr_data : cam_loc60;
	cam_loc61 <= (internal_wr_en & (internal_wr_ptr == 11'd61) ) ? wr_data : cam_loc61;
	cam_loc62 <= (internal_wr_en & (internal_wr_ptr == 11'd62) ) ? wr_data : cam_loc62;
	cam_loc63 <= (internal_wr_en & (internal_wr_ptr == 11'd63) ) ? wr_data : cam_loc63;
	cam_loc64 <= (internal_wr_en & (internal_wr_ptr == 11'd64) ) ? wr_data : cam_loc64;
	cam_loc65 <= (internal_wr_en & (internal_wr_ptr == 11'd65) ) ? wr_data : cam_loc65;
	cam_loc66 <= (internal_wr_en & (internal_wr_ptr == 11'd66) ) ? wr_data : cam_loc66;
	cam_loc67 <= (internal_wr_en & (internal_wr_ptr == 11'd67) ) ? wr_data : cam_loc67;
	cam_loc68 <= (internal_wr_en & (internal_wr_ptr == 11'd68) ) ? wr_data : cam_loc68;
	cam_loc69 <= (internal_wr_en & (internal_wr_ptr == 11'd69) ) ? wr_data : cam_loc69;
	cam_loc70 <= (internal_wr_en & (internal_wr_ptr == 11'd70) ) ? wr_data : cam_loc70;
	cam_loc71 <= (internal_wr_en & (internal_wr_ptr == 11'd71) ) ? wr_data : cam_loc71;
	cam_loc72 <= (internal_wr_en & (internal_wr_ptr == 11'd72) ) ? wr_data : cam_loc72;
	cam_loc73 <= (internal_wr_en & (internal_wr_ptr == 11'd73) ) ? wr_data : cam_loc73;
	cam_loc74 <= (internal_wr_en & (internal_wr_ptr == 11'd74) ) ? wr_data : cam_loc74;
	cam_loc75 <= (internal_wr_en & (internal_wr_ptr == 11'd75) ) ? wr_data : cam_loc75;
	cam_loc76 <= (internal_wr_en & (internal_wr_ptr == 11'd76) ) ? wr_data : cam_loc76;
	cam_loc77 <= (internal_wr_en & (internal_wr_ptr == 11'd77) ) ? wr_data : cam_loc77;
	cam_loc78 <= (internal_wr_en & (internal_wr_ptr == 11'd78) ) ? wr_data : cam_loc78;
	cam_loc79 <= (internal_wr_en & (internal_wr_ptr == 11'd79) ) ? wr_data : cam_loc79;
	cam_loc80 <= (internal_wr_en & (internal_wr_ptr == 11'd80) ) ? wr_data : cam_loc80;
	cam_loc81 <= (internal_wr_en & (internal_wr_ptr == 11'd81) ) ? wr_data : cam_loc81;
	cam_loc82 <= (internal_wr_en & (internal_wr_ptr == 11'd82) ) ? wr_data : cam_loc82;
	cam_loc83 <= (internal_wr_en & (internal_wr_ptr == 11'd83) ) ? wr_data : cam_loc83;
	cam_loc84 <= (internal_wr_en & (internal_wr_ptr == 11'd84) ) ? wr_data : cam_loc84;
	cam_loc85 <= (internal_wr_en & (internal_wr_ptr == 11'd85) ) ? wr_data : cam_loc85;
	cam_loc86 <= (internal_wr_en & (internal_wr_ptr == 11'd86) ) ? wr_data : cam_loc86;
	cam_loc87 <= (internal_wr_en & (internal_wr_ptr == 11'd87) ) ? wr_data : cam_loc87;
	cam_loc88 <= (internal_wr_en & (internal_wr_ptr == 11'd88) ) ? wr_data : cam_loc88;
	cam_loc89 <= (internal_wr_en & (internal_wr_ptr == 11'd89) ) ? wr_data : cam_loc89;
	cam_loc90 <= (internal_wr_en & (internal_wr_ptr == 11'd90) ) ? wr_data : cam_loc90;
	cam_loc91 <= (internal_wr_en & (internal_wr_ptr == 11'd91) ) ? wr_data : cam_loc91;
	cam_loc92 <= (internal_wr_en & (internal_wr_ptr == 11'd92) ) ? wr_data : cam_loc92;
	cam_loc93 <= (internal_wr_en & (internal_wr_ptr == 11'd93) ) ? wr_data : cam_loc93;
	cam_loc94 <= (internal_wr_en & (internal_wr_ptr == 11'd94) ) ? wr_data : cam_loc94;
	cam_loc95 <= (internal_wr_en & (internal_wr_ptr == 11'd95) ) ? wr_data : cam_loc95;
	cam_loc96 <= (internal_wr_en & (internal_wr_ptr == 11'd96) ) ? wr_data : cam_loc96;
	cam_loc97 <= (internal_wr_en & (internal_wr_ptr == 11'd97) ) ? wr_data : cam_loc97;
	cam_loc98 <= (internal_wr_en & (internal_wr_ptr == 11'd98) ) ? wr_data : cam_loc98;
	cam_loc99 <= (internal_wr_en & (internal_wr_ptr == 11'd99) ) ? wr_data : cam_loc99;
	cam_loc100 <= (internal_wr_en & (internal_wr_ptr == 11'd100) ) ? wr_data : cam_loc100;
	cam_loc101 <= (internal_wr_en & (internal_wr_ptr == 11'd101) ) ? wr_data : cam_loc101;
	cam_loc102 <= (internal_wr_en & (internal_wr_ptr == 11'd102) ) ? wr_data : cam_loc102;
	cam_loc103 <= (internal_wr_en & (internal_wr_ptr == 11'd103) ) ? wr_data : cam_loc103;
	cam_loc104 <= (internal_wr_en & (internal_wr_ptr == 11'd104) ) ? wr_data : cam_loc104;
	cam_loc105 <= (internal_wr_en & (internal_wr_ptr == 11'd105) ) ? wr_data : cam_loc105;
	cam_loc106 <= (internal_wr_en & (internal_wr_ptr == 11'd106) ) ? wr_data : cam_loc106;
	cam_loc107 <= (internal_wr_en & (internal_wr_ptr == 11'd107) ) ? wr_data : cam_loc107;
	cam_loc108 <= (internal_wr_en & (internal_wr_ptr == 11'd108) ) ? wr_data : cam_loc108;
	cam_loc109 <= (internal_wr_en & (internal_wr_ptr == 11'd109) ) ? wr_data : cam_loc109;
	cam_loc110 <= (internal_wr_en & (internal_wr_ptr == 11'd110) ) ? wr_data : cam_loc110;
	cam_loc111 <= (internal_wr_en & (internal_wr_ptr == 11'd111) ) ? wr_data : cam_loc111;
	cam_loc112 <= (internal_wr_en & (internal_wr_ptr == 11'd112) ) ? wr_data : cam_loc112;
	cam_loc113 <= (internal_wr_en & (internal_wr_ptr == 11'd113) ) ? wr_data : cam_loc113;
	cam_loc114 <= (internal_wr_en & (internal_wr_ptr == 11'd114) ) ? wr_data : cam_loc114;
	cam_loc115 <= (internal_wr_en & (internal_wr_ptr == 11'd115) ) ? wr_data : cam_loc115;
	cam_loc116 <= (internal_wr_en & (internal_wr_ptr == 11'd116) ) ? wr_data : cam_loc116;
	cam_loc117 <= (internal_wr_en & (internal_wr_ptr == 11'd117) ) ? wr_data : cam_loc117;
	cam_loc118 <= (internal_wr_en & (internal_wr_ptr == 11'd118) ) ? wr_data : cam_loc118;
	cam_loc119 <= (internal_wr_en & (internal_wr_ptr == 11'd119) ) ? wr_data : cam_loc119;
	cam_loc120 <= (internal_wr_en & (internal_wr_ptr == 11'd120) ) ? wr_data : cam_loc120;
	cam_loc121 <= (internal_wr_en & (internal_wr_ptr == 11'd121) ) ? wr_data : cam_loc121;
	cam_loc122 <= (internal_wr_en & (internal_wr_ptr == 11'd122) ) ? wr_data : cam_loc122;
	cam_loc123 <= (internal_wr_en & (internal_wr_ptr == 11'd123) ) ? wr_data : cam_loc123;
	cam_loc124 <= (internal_wr_en & (internal_wr_ptr == 11'd124) ) ? wr_data : cam_loc124;
	cam_loc125 <= (internal_wr_en & (internal_wr_ptr == 11'd125) ) ? wr_data : cam_loc125;
	cam_loc126 <= (internal_wr_en & (internal_wr_ptr == 11'd126) ) ? wr_data : cam_loc126;
	cam_loc127 <= (internal_wr_en & (internal_wr_ptr == 11'd127) ) ? wr_data : cam_loc127;
	cam_loc128 <= (internal_wr_en & (internal_wr_ptr == 11'd128) ) ? wr_data : cam_loc128;
	cam_loc129 <= (internal_wr_en & (internal_wr_ptr == 11'd129) ) ? wr_data : cam_loc129;
	cam_loc130 <= (internal_wr_en & (internal_wr_ptr == 11'd130) ) ? wr_data : cam_loc130;
	cam_loc131 <= (internal_wr_en & (internal_wr_ptr == 11'd131) ) ? wr_data : cam_loc131;
	cam_loc132 <= (internal_wr_en & (internal_wr_ptr == 11'd132) ) ? wr_data : cam_loc132;
	cam_loc133 <= (internal_wr_en & (internal_wr_ptr == 11'd133) ) ? wr_data : cam_loc133;
	cam_loc134 <= (internal_wr_en & (internal_wr_ptr == 11'd134) ) ? wr_data : cam_loc134;
	cam_loc135 <= (internal_wr_en & (internal_wr_ptr == 11'd135) ) ? wr_data : cam_loc135;
	cam_loc136 <= (internal_wr_en & (internal_wr_ptr == 11'd136) ) ? wr_data : cam_loc136;
	cam_loc137 <= (internal_wr_en & (internal_wr_ptr == 11'd137) ) ? wr_data : cam_loc137;
	cam_loc138 <= (internal_wr_en & (internal_wr_ptr == 11'd138) ) ? wr_data : cam_loc138;
	cam_loc139 <= (internal_wr_en & (internal_wr_ptr == 11'd139) ) ? wr_data : cam_loc139;
	cam_loc140 <= (internal_wr_en & (internal_wr_ptr == 11'd140) ) ? wr_data : cam_loc140;
	cam_loc141 <= (internal_wr_en & (internal_wr_ptr == 11'd141) ) ? wr_data : cam_loc141;
	cam_loc142 <= (internal_wr_en & (internal_wr_ptr == 11'd142) ) ? wr_data : cam_loc142;
	cam_loc143 <= (internal_wr_en & (internal_wr_ptr == 11'd143) ) ? wr_data : cam_loc143;
	cam_loc144 <= (internal_wr_en & (internal_wr_ptr == 11'd144) ) ? wr_data : cam_loc144;
	cam_loc145 <= (internal_wr_en & (internal_wr_ptr == 11'd145) ) ? wr_data : cam_loc145;
	cam_loc146 <= (internal_wr_en & (internal_wr_ptr == 11'd146) ) ? wr_data : cam_loc146;
	cam_loc147 <= (internal_wr_en & (internal_wr_ptr == 11'd147) ) ? wr_data : cam_loc147;
	cam_loc148 <= (internal_wr_en & (internal_wr_ptr == 11'd148) ) ? wr_data : cam_loc148;
	cam_loc149 <= (internal_wr_en & (internal_wr_ptr == 11'd149) ) ? wr_data : cam_loc149;
	cam_loc150 <= (internal_wr_en & (internal_wr_ptr == 11'd150) ) ? wr_data : cam_loc150;
	cam_loc151 <= (internal_wr_en & (internal_wr_ptr == 11'd151) ) ? wr_data : cam_loc151;
	cam_loc152 <= (internal_wr_en & (internal_wr_ptr == 11'd152) ) ? wr_data : cam_loc152;
	cam_loc153 <= (internal_wr_en & (internal_wr_ptr == 11'd153) ) ? wr_data : cam_loc153;
	cam_loc154 <= (internal_wr_en & (internal_wr_ptr == 11'd154) ) ? wr_data : cam_loc154;
	cam_loc155 <= (internal_wr_en & (internal_wr_ptr == 11'd155) ) ? wr_data : cam_loc155;
	cam_loc156 <= (internal_wr_en & (internal_wr_ptr == 11'd156) ) ? wr_data : cam_loc156;
	cam_loc157 <= (internal_wr_en & (internal_wr_ptr == 11'd157) ) ? wr_data : cam_loc157;
	cam_loc158 <= (internal_wr_en & (internal_wr_ptr == 11'd158) ) ? wr_data : cam_loc158;
	cam_loc159 <= (internal_wr_en & (internal_wr_ptr == 11'd159) ) ? wr_data : cam_loc159;
	cam_loc160 <= (internal_wr_en & (internal_wr_ptr == 11'd160) ) ? wr_data : cam_loc160;
	cam_loc161 <= (internal_wr_en & (internal_wr_ptr == 11'd161) ) ? wr_data : cam_loc161;
	cam_loc162 <= (internal_wr_en & (internal_wr_ptr == 11'd162) ) ? wr_data : cam_loc162;
	cam_loc163 <= (internal_wr_en & (internal_wr_ptr == 11'd163) ) ? wr_data : cam_loc163;
	cam_loc164 <= (internal_wr_en & (internal_wr_ptr == 11'd164) ) ? wr_data : cam_loc164;
	cam_loc165 <= (internal_wr_en & (internal_wr_ptr == 11'd165) ) ? wr_data : cam_loc165;
	cam_loc166 <= (internal_wr_en & (internal_wr_ptr == 11'd166) ) ? wr_data : cam_loc166;
	cam_loc167 <= (internal_wr_en & (internal_wr_ptr == 11'd167) ) ? wr_data : cam_loc167;
	cam_loc168 <= (internal_wr_en & (internal_wr_ptr == 11'd168) ) ? wr_data : cam_loc168;
	cam_loc169 <= (internal_wr_en & (internal_wr_ptr == 11'd169) ) ? wr_data : cam_loc169;
	cam_loc170 <= (internal_wr_en & (internal_wr_ptr == 11'd170) ) ? wr_data : cam_loc170;
	cam_loc171 <= (internal_wr_en & (internal_wr_ptr == 11'd171) ) ? wr_data : cam_loc171;
	cam_loc172 <= (internal_wr_en & (internal_wr_ptr == 11'd172) ) ? wr_data : cam_loc172;
	cam_loc173 <= (internal_wr_en & (internal_wr_ptr == 11'd173) ) ? wr_data : cam_loc173;
	cam_loc174 <= (internal_wr_en & (internal_wr_ptr == 11'd174) ) ? wr_data : cam_loc174;
	cam_loc175 <= (internal_wr_en & (internal_wr_ptr == 11'd175) ) ? wr_data : cam_loc175;
	cam_loc176 <= (internal_wr_en & (internal_wr_ptr == 11'd176) ) ? wr_data : cam_loc176;
	cam_loc177 <= (internal_wr_en & (internal_wr_ptr == 11'd177) ) ? wr_data : cam_loc177;
	cam_loc178 <= (internal_wr_en & (internal_wr_ptr == 11'd178) ) ? wr_data : cam_loc178;
	cam_loc179 <= (internal_wr_en & (internal_wr_ptr == 11'd179) ) ? wr_data : cam_loc179;
	cam_loc180 <= (internal_wr_en & (internal_wr_ptr == 11'd180) ) ? wr_data : cam_loc180;
	cam_loc181 <= (internal_wr_en & (internal_wr_ptr == 11'd181) ) ? wr_data : cam_loc181;
	cam_loc182 <= (internal_wr_en & (internal_wr_ptr == 11'd182) ) ? wr_data : cam_loc182;
	cam_loc183 <= (internal_wr_en & (internal_wr_ptr == 11'd183) ) ? wr_data : cam_loc183;
	cam_loc184 <= (internal_wr_en & (internal_wr_ptr == 11'd184) ) ? wr_data : cam_loc184;
	cam_loc185 <= (internal_wr_en & (internal_wr_ptr == 11'd185) ) ? wr_data : cam_loc185;
	cam_loc186 <= (internal_wr_en & (internal_wr_ptr == 11'd186) ) ? wr_data : cam_loc186;
	cam_loc187 <= (internal_wr_en & (internal_wr_ptr == 11'd187) ) ? wr_data : cam_loc187;
	cam_loc188 <= (internal_wr_en & (internal_wr_ptr == 11'd188) ) ? wr_data : cam_loc188;
	cam_loc189 <= (internal_wr_en & (internal_wr_ptr == 11'd189) ) ? wr_data : cam_loc189;
	cam_loc190 <= (internal_wr_en & (internal_wr_ptr == 11'd190) ) ? wr_data : cam_loc190;
	cam_loc191 <= (internal_wr_en & (internal_wr_ptr == 11'd191) ) ? wr_data : cam_loc191;
	cam_loc192 <= (internal_wr_en & (internal_wr_ptr == 11'd192) ) ? wr_data : cam_loc192;
	cam_loc193 <= (internal_wr_en & (internal_wr_ptr == 11'd193) ) ? wr_data : cam_loc193;
	cam_loc194 <= (internal_wr_en & (internal_wr_ptr == 11'd194) ) ? wr_data : cam_loc194;
	cam_loc195 <= (internal_wr_en & (internal_wr_ptr == 11'd195) ) ? wr_data : cam_loc195;
	cam_loc196 <= (internal_wr_en & (internal_wr_ptr == 11'd196) ) ? wr_data : cam_loc196;
	cam_loc197 <= (internal_wr_en & (internal_wr_ptr == 11'd197) ) ? wr_data : cam_loc197;
	cam_loc198 <= (internal_wr_en & (internal_wr_ptr == 11'd198) ) ? wr_data : cam_loc198;
	cam_loc199 <= (internal_wr_en & (internal_wr_ptr == 11'd199) ) ? wr_data : cam_loc199;
	cam_loc200 <= (internal_wr_en & (internal_wr_ptr == 11'd200) ) ? wr_data : cam_loc200;
	cam_loc201 <= (internal_wr_en & (internal_wr_ptr == 11'd201) ) ? wr_data : cam_loc201;
	cam_loc202 <= (internal_wr_en & (internal_wr_ptr == 11'd202) ) ? wr_data : cam_loc202;
	cam_loc203 <= (internal_wr_en & (internal_wr_ptr == 11'd203) ) ? wr_data : cam_loc203;
	cam_loc204 <= (internal_wr_en & (internal_wr_ptr == 11'd204) ) ? wr_data : cam_loc204;
	cam_loc205 <= (internal_wr_en & (internal_wr_ptr == 11'd205) ) ? wr_data : cam_loc205;
	cam_loc206 <= (internal_wr_en & (internal_wr_ptr == 11'd206) ) ? wr_data : cam_loc206;
	cam_loc207 <= (internal_wr_en & (internal_wr_ptr == 11'd207) ) ? wr_data : cam_loc207;
	cam_loc208 <= (internal_wr_en & (internal_wr_ptr == 11'd208) ) ? wr_data : cam_loc208;
	cam_loc209 <= (internal_wr_en & (internal_wr_ptr == 11'd209) ) ? wr_data : cam_loc209;
	cam_loc210 <= (internal_wr_en & (internal_wr_ptr == 11'd210) ) ? wr_data : cam_loc210;
	cam_loc211 <= (internal_wr_en & (internal_wr_ptr == 11'd211) ) ? wr_data : cam_loc211;
	cam_loc212 <= (internal_wr_en & (internal_wr_ptr == 11'd212) ) ? wr_data : cam_loc212;
	cam_loc213 <= (internal_wr_en & (internal_wr_ptr == 11'd213) ) ? wr_data : cam_loc213;
	cam_loc214 <= (internal_wr_en & (internal_wr_ptr == 11'd214) ) ? wr_data : cam_loc214;
	cam_loc215 <= (internal_wr_en & (internal_wr_ptr == 11'd215) ) ? wr_data : cam_loc215;
	cam_loc216 <= (internal_wr_en & (internal_wr_ptr == 11'd216) ) ? wr_data : cam_loc216;
	cam_loc217 <= (internal_wr_en & (internal_wr_ptr == 11'd217) ) ? wr_data : cam_loc217;
	cam_loc218 <= (internal_wr_en & (internal_wr_ptr == 11'd218) ) ? wr_data : cam_loc218;
	cam_loc219 <= (internal_wr_en & (internal_wr_ptr == 11'd219) ) ? wr_data : cam_loc219;
	cam_loc220 <= (internal_wr_en & (internal_wr_ptr == 11'd220) ) ? wr_data : cam_loc220;
	cam_loc221 <= (internal_wr_en & (internal_wr_ptr == 11'd221) ) ? wr_data : cam_loc221;
	cam_loc222 <= (internal_wr_en & (internal_wr_ptr == 11'd222) ) ? wr_data : cam_loc222;
	cam_loc223 <= (internal_wr_en & (internal_wr_ptr == 11'd223) ) ? wr_data : cam_loc223;
	cam_loc224 <= (internal_wr_en & (internal_wr_ptr == 11'd224) ) ? wr_data : cam_loc224;
	cam_loc225 <= (internal_wr_en & (internal_wr_ptr == 11'd225) ) ? wr_data : cam_loc225;
	cam_loc226 <= (internal_wr_en & (internal_wr_ptr == 11'd226) ) ? wr_data : cam_loc226;
	cam_loc227 <= (internal_wr_en & (internal_wr_ptr == 11'd227) ) ? wr_data : cam_loc227;
	cam_loc228 <= (internal_wr_en & (internal_wr_ptr == 11'd228) ) ? wr_data : cam_loc228;
	cam_loc229 <= (internal_wr_en & (internal_wr_ptr == 11'd229) ) ? wr_data : cam_loc229;
	cam_loc230 <= (internal_wr_en & (internal_wr_ptr == 11'd230) ) ? wr_data : cam_loc230;
	cam_loc231 <= (internal_wr_en & (internal_wr_ptr == 11'd231) ) ? wr_data : cam_loc231;
	cam_loc232 <= (internal_wr_en & (internal_wr_ptr == 11'd232) ) ? wr_data : cam_loc232;
	cam_loc233 <= (internal_wr_en & (internal_wr_ptr == 11'd233) ) ? wr_data : cam_loc233;
	cam_loc234 <= (internal_wr_en & (internal_wr_ptr == 11'd234) ) ? wr_data : cam_loc234;
	cam_loc235 <= (internal_wr_en & (internal_wr_ptr == 11'd235) ) ? wr_data : cam_loc235;
	cam_loc236 <= (internal_wr_en & (internal_wr_ptr == 11'd236) ) ? wr_data : cam_loc236;
	cam_loc237 <= (internal_wr_en & (internal_wr_ptr == 11'd237) ) ? wr_data : cam_loc237;
	cam_loc238 <= (internal_wr_en & (internal_wr_ptr == 11'd238) ) ? wr_data : cam_loc238;
	cam_loc239 <= (internal_wr_en & (internal_wr_ptr == 11'd239) ) ? wr_data : cam_loc239;
	cam_loc240 <= (internal_wr_en & (internal_wr_ptr == 11'd240) ) ? wr_data : cam_loc240;
	cam_loc241 <= (internal_wr_en & (internal_wr_ptr == 11'd241) ) ? wr_data : cam_loc241;
	cam_loc242 <= (internal_wr_en & (internal_wr_ptr == 11'd242) ) ? wr_data : cam_loc242;
	cam_loc243 <= (internal_wr_en & (internal_wr_ptr == 11'd243) ) ? wr_data : cam_loc243;
	cam_loc244 <= (internal_wr_en & (internal_wr_ptr == 11'd244) ) ? wr_data : cam_loc244;
	cam_loc245 <= (internal_wr_en & (internal_wr_ptr == 11'd245) ) ? wr_data : cam_loc245;
	cam_loc246 <= (internal_wr_en & (internal_wr_ptr == 11'd246) ) ? wr_data : cam_loc246;
	cam_loc247 <= (internal_wr_en & (internal_wr_ptr == 11'd247) ) ? wr_data : cam_loc247;
	cam_loc248 <= (internal_wr_en & (internal_wr_ptr == 11'd248) ) ? wr_data : cam_loc248;
	cam_loc249 <= (internal_wr_en & (internal_wr_ptr == 11'd249) ) ? wr_data : cam_loc249;
	cam_loc250 <= (internal_wr_en & (internal_wr_ptr == 11'd250) ) ? wr_data : cam_loc250;
	cam_loc251 <= (internal_wr_en & (internal_wr_ptr == 11'd251) ) ? wr_data : cam_loc251;
	cam_loc252 <= (internal_wr_en & (internal_wr_ptr == 11'd252) ) ? wr_data : cam_loc252;
	cam_loc253 <= (internal_wr_en & (internal_wr_ptr == 11'd253) ) ? wr_data : cam_loc253;
	cam_loc254 <= (internal_wr_en & (internal_wr_ptr == 11'd254) ) ? wr_data : cam_loc254;
	cam_loc255 <= (internal_wr_en & (internal_wr_ptr == 11'd255) ) ? wr_data : cam_loc255;
	cam_loc256 <= (internal_wr_en & (internal_wr_ptr == 11'd256) ) ? wr_data : cam_loc256;
	cam_loc257 <= (internal_wr_en & (internal_wr_ptr == 11'd257) ) ? wr_data : cam_loc257;
	cam_loc258 <= (internal_wr_en & (internal_wr_ptr == 11'd258) ) ? wr_data : cam_loc258;
	cam_loc259 <= (internal_wr_en & (internal_wr_ptr == 11'd259) ) ? wr_data : cam_loc259;
	cam_loc260 <= (internal_wr_en & (internal_wr_ptr == 11'd260) ) ? wr_data : cam_loc260;
	cam_loc261 <= (internal_wr_en & (internal_wr_ptr == 11'd261) ) ? wr_data : cam_loc261;
	cam_loc262 <= (internal_wr_en & (internal_wr_ptr == 11'd262) ) ? wr_data : cam_loc262;
	cam_loc263 <= (internal_wr_en & (internal_wr_ptr == 11'd263) ) ? wr_data : cam_loc263;
	cam_loc264 <= (internal_wr_en & (internal_wr_ptr == 11'd264) ) ? wr_data : cam_loc264;
	cam_loc265 <= (internal_wr_en & (internal_wr_ptr == 11'd265) ) ? wr_data : cam_loc265;
	cam_loc266 <= (internal_wr_en & (internal_wr_ptr == 11'd266) ) ? wr_data : cam_loc266;
	cam_loc267 <= (internal_wr_en & (internal_wr_ptr == 11'd267) ) ? wr_data : cam_loc267;
	cam_loc268 <= (internal_wr_en & (internal_wr_ptr == 11'd268) ) ? wr_data : cam_loc268;
	cam_loc269 <= (internal_wr_en & (internal_wr_ptr == 11'd269) ) ? wr_data : cam_loc269;
	cam_loc270 <= (internal_wr_en & (internal_wr_ptr == 11'd270) ) ? wr_data : cam_loc270;
	cam_loc271 <= (internal_wr_en & (internal_wr_ptr == 11'd271) ) ? wr_data : cam_loc271;
	cam_loc272 <= (internal_wr_en & (internal_wr_ptr == 11'd272) ) ? wr_data : cam_loc272;
	cam_loc273 <= (internal_wr_en & (internal_wr_ptr == 11'd273) ) ? wr_data : cam_loc273;
	cam_loc274 <= (internal_wr_en & (internal_wr_ptr == 11'd274) ) ? wr_data : cam_loc274;
	cam_loc275 <= (internal_wr_en & (internal_wr_ptr == 11'd275) ) ? wr_data : cam_loc275;
	cam_loc276 <= (internal_wr_en & (internal_wr_ptr == 11'd276) ) ? wr_data : cam_loc276;
	cam_loc277 <= (internal_wr_en & (internal_wr_ptr == 11'd277) ) ? wr_data : cam_loc277;
	cam_loc278 <= (internal_wr_en & (internal_wr_ptr == 11'd278) ) ? wr_data : cam_loc278;
	cam_loc279 <= (internal_wr_en & (internal_wr_ptr == 11'd279) ) ? wr_data : cam_loc279;
	cam_loc280 <= (internal_wr_en & (internal_wr_ptr == 11'd280) ) ? wr_data : cam_loc280;
	cam_loc281 <= (internal_wr_en & (internal_wr_ptr == 11'd281) ) ? wr_data : cam_loc281;
	cam_loc282 <= (internal_wr_en & (internal_wr_ptr == 11'd282) ) ? wr_data : cam_loc282;
	cam_loc283 <= (internal_wr_en & (internal_wr_ptr == 11'd283) ) ? wr_data : cam_loc283;
	cam_loc284 <= (internal_wr_en & (internal_wr_ptr == 11'd284) ) ? wr_data : cam_loc284;
	cam_loc285 <= (internal_wr_en & (internal_wr_ptr == 11'd285) ) ? wr_data : cam_loc285;
	cam_loc286 <= (internal_wr_en & (internal_wr_ptr == 11'd286) ) ? wr_data : cam_loc286;
	cam_loc287 <= (internal_wr_en & (internal_wr_ptr == 11'd287) ) ? wr_data : cam_loc287;
	cam_loc288 <= (internal_wr_en & (internal_wr_ptr == 11'd288) ) ? wr_data : cam_loc288;
	cam_loc289 <= (internal_wr_en & (internal_wr_ptr == 11'd289) ) ? wr_data : cam_loc289;
	cam_loc290 <= (internal_wr_en & (internal_wr_ptr == 11'd290) ) ? wr_data : cam_loc290;
	cam_loc291 <= (internal_wr_en & (internal_wr_ptr == 11'd291) ) ? wr_data : cam_loc291;
	cam_loc292 <= (internal_wr_en & (internal_wr_ptr == 11'd292) ) ? wr_data : cam_loc292;
	cam_loc293 <= (internal_wr_en & (internal_wr_ptr == 11'd293) ) ? wr_data : cam_loc293;
	cam_loc294 <= (internal_wr_en & (internal_wr_ptr == 11'd294) ) ? wr_data : cam_loc294;
	cam_loc295 <= (internal_wr_en & (internal_wr_ptr == 11'd295) ) ? wr_data : cam_loc295;
	cam_loc296 <= (internal_wr_en & (internal_wr_ptr == 11'd296) ) ? wr_data : cam_loc296;
	cam_loc297 <= (internal_wr_en & (internal_wr_ptr == 11'd297) ) ? wr_data : cam_loc297;
	cam_loc298 <= (internal_wr_en & (internal_wr_ptr == 11'd298) ) ? wr_data : cam_loc298;
	cam_loc299 <= (internal_wr_en & (internal_wr_ptr == 11'd299) ) ? wr_data : cam_loc299;
	cam_loc300 <= (internal_wr_en & (internal_wr_ptr == 11'd300) ) ? wr_data : cam_loc300;
	cam_loc301 <= (internal_wr_en & (internal_wr_ptr == 11'd301) ) ? wr_data : cam_loc301;
	cam_loc302 <= (internal_wr_en & (internal_wr_ptr == 11'd302) ) ? wr_data : cam_loc302;
	cam_loc303 <= (internal_wr_en & (internal_wr_ptr == 11'd303) ) ? wr_data : cam_loc303;
	cam_loc304 <= (internal_wr_en & (internal_wr_ptr == 11'd304) ) ? wr_data : cam_loc304;
	cam_loc305 <= (internal_wr_en & (internal_wr_ptr == 11'd305) ) ? wr_data : cam_loc305;
	cam_loc306 <= (internal_wr_en & (internal_wr_ptr == 11'd306) ) ? wr_data : cam_loc306;
	cam_loc307 <= (internal_wr_en & (internal_wr_ptr == 11'd307) ) ? wr_data : cam_loc307;
	cam_loc308 <= (internal_wr_en & (internal_wr_ptr == 11'd308) ) ? wr_data : cam_loc308;
	cam_loc309 <= (internal_wr_en & (internal_wr_ptr == 11'd309) ) ? wr_data : cam_loc309;
	cam_loc310 <= (internal_wr_en & (internal_wr_ptr == 11'd310) ) ? wr_data : cam_loc310;
	cam_loc311 <= (internal_wr_en & (internal_wr_ptr == 11'd311) ) ? wr_data : cam_loc311;
	cam_loc312 <= (internal_wr_en & (internal_wr_ptr == 11'd312) ) ? wr_data : cam_loc312;
	cam_loc313 <= (internal_wr_en & (internal_wr_ptr == 11'd313) ) ? wr_data : cam_loc313;
	cam_loc314 <= (internal_wr_en & (internal_wr_ptr == 11'd314) ) ? wr_data : cam_loc314;
	cam_loc315 <= (internal_wr_en & (internal_wr_ptr == 11'd315) ) ? wr_data : cam_loc315;
	cam_loc316 <= (internal_wr_en & (internal_wr_ptr == 11'd316) ) ? wr_data : cam_loc316;
	cam_loc317 <= (internal_wr_en & (internal_wr_ptr == 11'd317) ) ? wr_data : cam_loc317;
	cam_loc318 <= (internal_wr_en & (internal_wr_ptr == 11'd318) ) ? wr_data : cam_loc318;
	cam_loc319 <= (internal_wr_en & (internal_wr_ptr == 11'd319) ) ? wr_data : cam_loc319;
	cam_loc320 <= (internal_wr_en & (internal_wr_ptr == 11'd320) ) ? wr_data : cam_loc320;
	cam_loc321 <= (internal_wr_en & (internal_wr_ptr == 11'd321) ) ? wr_data : cam_loc321;
	cam_loc322 <= (internal_wr_en & (internal_wr_ptr == 11'd322) ) ? wr_data : cam_loc322;
	cam_loc323 <= (internal_wr_en & (internal_wr_ptr == 11'd323) ) ? wr_data : cam_loc323;
	cam_loc324 <= (internal_wr_en & (internal_wr_ptr == 11'd324) ) ? wr_data : cam_loc324;
	cam_loc325 <= (internal_wr_en & (internal_wr_ptr == 11'd325) ) ? wr_data : cam_loc325;
	cam_loc326 <= (internal_wr_en & (internal_wr_ptr == 11'd326) ) ? wr_data : cam_loc326;
	cam_loc327 <= (internal_wr_en & (internal_wr_ptr == 11'd327) ) ? wr_data : cam_loc327;
	cam_loc328 <= (internal_wr_en & (internal_wr_ptr == 11'd328) ) ? wr_data : cam_loc328;
	cam_loc329 <= (internal_wr_en & (internal_wr_ptr == 11'd329) ) ? wr_data : cam_loc329;
	cam_loc330 <= (internal_wr_en & (internal_wr_ptr == 11'd330) ) ? wr_data : cam_loc330;
	cam_loc331 <= (internal_wr_en & (internal_wr_ptr == 11'd331) ) ? wr_data : cam_loc331;
	cam_loc332 <= (internal_wr_en & (internal_wr_ptr == 11'd332) ) ? wr_data : cam_loc332;
	cam_loc333 <= (internal_wr_en & (internal_wr_ptr == 11'd333) ) ? wr_data : cam_loc333;
	cam_loc334 <= (internal_wr_en & (internal_wr_ptr == 11'd334) ) ? wr_data : cam_loc334;
	cam_loc335 <= (internal_wr_en & (internal_wr_ptr == 11'd335) ) ? wr_data : cam_loc335;
	cam_loc336 <= (internal_wr_en & (internal_wr_ptr == 11'd336) ) ? wr_data : cam_loc336;
	cam_loc337 <= (internal_wr_en & (internal_wr_ptr == 11'd337) ) ? wr_data : cam_loc337;
	cam_loc338 <= (internal_wr_en & (internal_wr_ptr == 11'd338) ) ? wr_data : cam_loc338;
	cam_loc339 <= (internal_wr_en & (internal_wr_ptr == 11'd339) ) ? wr_data : cam_loc339;
	cam_loc340 <= (internal_wr_en & (internal_wr_ptr == 11'd340) ) ? wr_data : cam_loc340;
	cam_loc341 <= (internal_wr_en & (internal_wr_ptr == 11'd341) ) ? wr_data : cam_loc341;
	cam_loc342 <= (internal_wr_en & (internal_wr_ptr == 11'd342) ) ? wr_data : cam_loc342;
	cam_loc343 <= (internal_wr_en & (internal_wr_ptr == 11'd343) ) ? wr_data : cam_loc343;
	cam_loc344 <= (internal_wr_en & (internal_wr_ptr == 11'd344) ) ? wr_data : cam_loc344;
	cam_loc345 <= (internal_wr_en & (internal_wr_ptr == 11'd345) ) ? wr_data : cam_loc345;
	cam_loc346 <= (internal_wr_en & (internal_wr_ptr == 11'd346) ) ? wr_data : cam_loc346;
	cam_loc347 <= (internal_wr_en & (internal_wr_ptr == 11'd347) ) ? wr_data : cam_loc347;
	cam_loc348 <= (internal_wr_en & (internal_wr_ptr == 11'd348) ) ? wr_data : cam_loc348;
	cam_loc349 <= (internal_wr_en & (internal_wr_ptr == 11'd349) ) ? wr_data : cam_loc349;
	cam_loc350 <= (internal_wr_en & (internal_wr_ptr == 11'd350) ) ? wr_data : cam_loc350;
	cam_loc351 <= (internal_wr_en & (internal_wr_ptr == 11'd351) ) ? wr_data : cam_loc351;
	cam_loc352 <= (internal_wr_en & (internal_wr_ptr == 11'd352) ) ? wr_data : cam_loc352;
	cam_loc353 <= (internal_wr_en & (internal_wr_ptr == 11'd353) ) ? wr_data : cam_loc353;
	cam_loc354 <= (internal_wr_en & (internal_wr_ptr == 11'd354) ) ? wr_data : cam_loc354;
	cam_loc355 <= (internal_wr_en & (internal_wr_ptr == 11'd355) ) ? wr_data : cam_loc355;
	cam_loc356 <= (internal_wr_en & (internal_wr_ptr == 11'd356) ) ? wr_data : cam_loc356;
	cam_loc357 <= (internal_wr_en & (internal_wr_ptr == 11'd357) ) ? wr_data : cam_loc357;
	cam_loc358 <= (internal_wr_en & (internal_wr_ptr == 11'd358) ) ? wr_data : cam_loc358;
	cam_loc359 <= (internal_wr_en & (internal_wr_ptr == 11'd359) ) ? wr_data : cam_loc359;
	cam_loc360 <= (internal_wr_en & (internal_wr_ptr == 11'd360) ) ? wr_data : cam_loc360;
	cam_loc361 <= (internal_wr_en & (internal_wr_ptr == 11'd361) ) ? wr_data : cam_loc361;
	cam_loc362 <= (internal_wr_en & (internal_wr_ptr == 11'd362) ) ? wr_data : cam_loc362;
	cam_loc363 <= (internal_wr_en & (internal_wr_ptr == 11'd363) ) ? wr_data : cam_loc363;
	cam_loc364 <= (internal_wr_en & (internal_wr_ptr == 11'd364) ) ? wr_data : cam_loc364;
	cam_loc365 <= (internal_wr_en & (internal_wr_ptr == 11'd365) ) ? wr_data : cam_loc365;
	cam_loc366 <= (internal_wr_en & (internal_wr_ptr == 11'd366) ) ? wr_data : cam_loc366;
	cam_loc367 <= (internal_wr_en & (internal_wr_ptr == 11'd367) ) ? wr_data : cam_loc367;
	cam_loc368 <= (internal_wr_en & (internal_wr_ptr == 11'd368) ) ? wr_data : cam_loc368;
	cam_loc369 <= (internal_wr_en & (internal_wr_ptr == 11'd369) ) ? wr_data : cam_loc369;
	cam_loc370 <= (internal_wr_en & (internal_wr_ptr == 11'd370) ) ? wr_data : cam_loc370;
	cam_loc371 <= (internal_wr_en & (internal_wr_ptr == 11'd371) ) ? wr_data : cam_loc371;
	cam_loc372 <= (internal_wr_en & (internal_wr_ptr == 11'd372) ) ? wr_data : cam_loc372;
	cam_loc373 <= (internal_wr_en & (internal_wr_ptr == 11'd373) ) ? wr_data : cam_loc373;
	cam_loc374 <= (internal_wr_en & (internal_wr_ptr == 11'd374) ) ? wr_data : cam_loc374;
	cam_loc375 <= (internal_wr_en & (internal_wr_ptr == 11'd375) ) ? wr_data : cam_loc375;
	cam_loc376 <= (internal_wr_en & (internal_wr_ptr == 11'd376) ) ? wr_data : cam_loc376;
	cam_loc377 <= (internal_wr_en & (internal_wr_ptr == 11'd377) ) ? wr_data : cam_loc377;
	cam_loc378 <= (internal_wr_en & (internal_wr_ptr == 11'd378) ) ? wr_data : cam_loc378;
	cam_loc379 <= (internal_wr_en & (internal_wr_ptr == 11'd379) ) ? wr_data : cam_loc379;
	cam_loc380 <= (internal_wr_en & (internal_wr_ptr == 11'd380) ) ? wr_data : cam_loc380;
	cam_loc381 <= (internal_wr_en & (internal_wr_ptr == 11'd381) ) ? wr_data : cam_loc381;
	cam_loc382 <= (internal_wr_en & (internal_wr_ptr == 11'd382) ) ? wr_data : cam_loc382;
	cam_loc383 <= (internal_wr_en & (internal_wr_ptr == 11'd383) ) ? wr_data : cam_loc383;
	cam_loc384 <= (internal_wr_en & (internal_wr_ptr == 11'd384) ) ? wr_data : cam_loc384;
	cam_loc385 <= (internal_wr_en & (internal_wr_ptr == 11'd385) ) ? wr_data : cam_loc385;
	cam_loc386 <= (internal_wr_en & (internal_wr_ptr == 11'd386) ) ? wr_data : cam_loc386;
	cam_loc387 <= (internal_wr_en & (internal_wr_ptr == 11'd387) ) ? wr_data : cam_loc387;
	cam_loc388 <= (internal_wr_en & (internal_wr_ptr == 11'd388) ) ? wr_data : cam_loc388;
	cam_loc389 <= (internal_wr_en & (internal_wr_ptr == 11'd389) ) ? wr_data : cam_loc389;
	cam_loc390 <= (internal_wr_en & (internal_wr_ptr == 11'd390) ) ? wr_data : cam_loc390;
	cam_loc391 <= (internal_wr_en & (internal_wr_ptr == 11'd391) ) ? wr_data : cam_loc391;
	cam_loc392 <= (internal_wr_en & (internal_wr_ptr == 11'd392) ) ? wr_data : cam_loc392;
	cam_loc393 <= (internal_wr_en & (internal_wr_ptr == 11'd393) ) ? wr_data : cam_loc393;
	cam_loc394 <= (internal_wr_en & (internal_wr_ptr == 11'd394) ) ? wr_data : cam_loc394;
	cam_loc395 <= (internal_wr_en & (internal_wr_ptr == 11'd395) ) ? wr_data : cam_loc395;
	cam_loc396 <= (internal_wr_en & (internal_wr_ptr == 11'd396) ) ? wr_data : cam_loc396;
	cam_loc397 <= (internal_wr_en & (internal_wr_ptr == 11'd397) ) ? wr_data : cam_loc397;
	cam_loc398 <= (internal_wr_en & (internal_wr_ptr == 11'd398) ) ? wr_data : cam_loc398;
	cam_loc399 <= (internal_wr_en & (internal_wr_ptr == 11'd399) ) ? wr_data : cam_loc399;
	cam_loc400 <= (internal_wr_en & (internal_wr_ptr == 11'd400) ) ? wr_data : cam_loc400;
	cam_loc401 <= (internal_wr_en & (internal_wr_ptr == 11'd401) ) ? wr_data : cam_loc401;
	cam_loc402 <= (internal_wr_en & (internal_wr_ptr == 11'd402) ) ? wr_data : cam_loc402;
	cam_loc403 <= (internal_wr_en & (internal_wr_ptr == 11'd403) ) ? wr_data : cam_loc403;
	cam_loc404 <= (internal_wr_en & (internal_wr_ptr == 11'd404) ) ? wr_data : cam_loc404;
	cam_loc405 <= (internal_wr_en & (internal_wr_ptr == 11'd405) ) ? wr_data : cam_loc405;
	cam_loc406 <= (internal_wr_en & (internal_wr_ptr == 11'd406) ) ? wr_data : cam_loc406;
	cam_loc407 <= (internal_wr_en & (internal_wr_ptr == 11'd407) ) ? wr_data : cam_loc407;
	cam_loc408 <= (internal_wr_en & (internal_wr_ptr == 11'd408) ) ? wr_data : cam_loc408;
	cam_loc409 <= (internal_wr_en & (internal_wr_ptr == 11'd409) ) ? wr_data : cam_loc409;
	cam_loc410 <= (internal_wr_en & (internal_wr_ptr == 11'd410) ) ? wr_data : cam_loc410;
	cam_loc411 <= (internal_wr_en & (internal_wr_ptr == 11'd411) ) ? wr_data : cam_loc411;
	cam_loc412 <= (internal_wr_en & (internal_wr_ptr == 11'd412) ) ? wr_data : cam_loc412;
	cam_loc413 <= (internal_wr_en & (internal_wr_ptr == 11'd413) ) ? wr_data : cam_loc413;
	cam_loc414 <= (internal_wr_en & (internal_wr_ptr == 11'd414) ) ? wr_data : cam_loc414;
	cam_loc415 <= (internal_wr_en & (internal_wr_ptr == 11'd415) ) ? wr_data : cam_loc415;
	cam_loc416 <= (internal_wr_en & (internal_wr_ptr == 11'd416) ) ? wr_data : cam_loc416;
	cam_loc417 <= (internal_wr_en & (internal_wr_ptr == 11'd417) ) ? wr_data : cam_loc417;
	cam_loc418 <= (internal_wr_en & (internal_wr_ptr == 11'd418) ) ? wr_data : cam_loc418;
	cam_loc419 <= (internal_wr_en & (internal_wr_ptr == 11'd419) ) ? wr_data : cam_loc419;
	cam_loc420 <= (internal_wr_en & (internal_wr_ptr == 11'd420) ) ? wr_data : cam_loc420;
	cam_loc421 <= (internal_wr_en & (internal_wr_ptr == 11'd421) ) ? wr_data : cam_loc421;
	cam_loc422 <= (internal_wr_en & (internal_wr_ptr == 11'd422) ) ? wr_data : cam_loc422;
	cam_loc423 <= (internal_wr_en & (internal_wr_ptr == 11'd423) ) ? wr_data : cam_loc423;
	cam_loc424 <= (internal_wr_en & (internal_wr_ptr == 11'd424) ) ? wr_data : cam_loc424;
	cam_loc425 <= (internal_wr_en & (internal_wr_ptr == 11'd425) ) ? wr_data : cam_loc425;
	cam_loc426 <= (internal_wr_en & (internal_wr_ptr == 11'd426) ) ? wr_data : cam_loc426;
	cam_loc427 <= (internal_wr_en & (internal_wr_ptr == 11'd427) ) ? wr_data : cam_loc427;
	cam_loc428 <= (internal_wr_en & (internal_wr_ptr == 11'd428) ) ? wr_data : cam_loc428;
	cam_loc429 <= (internal_wr_en & (internal_wr_ptr == 11'd429) ) ? wr_data : cam_loc429;
	cam_loc430 <= (internal_wr_en & (internal_wr_ptr == 11'd430) ) ? wr_data : cam_loc430;
	cam_loc431 <= (internal_wr_en & (internal_wr_ptr == 11'd431) ) ? wr_data : cam_loc431;
	cam_loc432 <= (internal_wr_en & (internal_wr_ptr == 11'd432) ) ? wr_data : cam_loc432;
	cam_loc433 <= (internal_wr_en & (internal_wr_ptr == 11'd433) ) ? wr_data : cam_loc433;
	cam_loc434 <= (internal_wr_en & (internal_wr_ptr == 11'd434) ) ? wr_data : cam_loc434;
	cam_loc435 <= (internal_wr_en & (internal_wr_ptr == 11'd435) ) ? wr_data : cam_loc435;
	cam_loc436 <= (internal_wr_en & (internal_wr_ptr == 11'd436) ) ? wr_data : cam_loc436;
	cam_loc437 <= (internal_wr_en & (internal_wr_ptr == 11'd437) ) ? wr_data : cam_loc437;
	cam_loc438 <= (internal_wr_en & (internal_wr_ptr == 11'd438) ) ? wr_data : cam_loc438;
	cam_loc439 <= (internal_wr_en & (internal_wr_ptr == 11'd439) ) ? wr_data : cam_loc439;
	cam_loc440 <= (internal_wr_en & (internal_wr_ptr == 11'd440) ) ? wr_data : cam_loc440;
	cam_loc441 <= (internal_wr_en & (internal_wr_ptr == 11'd441) ) ? wr_data : cam_loc441;
	cam_loc442 <= (internal_wr_en & (internal_wr_ptr == 11'd442) ) ? wr_data : cam_loc442;
	cam_loc443 <= (internal_wr_en & (internal_wr_ptr == 11'd443) ) ? wr_data : cam_loc443;
	cam_loc444 <= (internal_wr_en & (internal_wr_ptr == 11'd444) ) ? wr_data : cam_loc444;
	cam_loc445 <= (internal_wr_en & (internal_wr_ptr == 11'd445) ) ? wr_data : cam_loc445;
	cam_loc446 <= (internal_wr_en & (internal_wr_ptr == 11'd446) ) ? wr_data : cam_loc446;
	cam_loc447 <= (internal_wr_en & (internal_wr_ptr == 11'd447) ) ? wr_data : cam_loc447;
	cam_loc448 <= (internal_wr_en & (internal_wr_ptr == 11'd448) ) ? wr_data : cam_loc448;
	cam_loc449 <= (internal_wr_en & (internal_wr_ptr == 11'd449) ) ? wr_data : cam_loc449;
	cam_loc450 <= (internal_wr_en & (internal_wr_ptr == 11'd450) ) ? wr_data : cam_loc450;
	cam_loc451 <= (internal_wr_en & (internal_wr_ptr == 11'd451) ) ? wr_data : cam_loc451;
	cam_loc452 <= (internal_wr_en & (internal_wr_ptr == 11'd452) ) ? wr_data : cam_loc452;
	cam_loc453 <= (internal_wr_en & (internal_wr_ptr == 11'd453) ) ? wr_data : cam_loc453;
	cam_loc454 <= (internal_wr_en & (internal_wr_ptr == 11'd454) ) ? wr_data : cam_loc454;
	cam_loc455 <= (internal_wr_en & (internal_wr_ptr == 11'd455) ) ? wr_data : cam_loc455;
	cam_loc456 <= (internal_wr_en & (internal_wr_ptr == 11'd456) ) ? wr_data : cam_loc456;
	cam_loc457 <= (internal_wr_en & (internal_wr_ptr == 11'd457) ) ? wr_data : cam_loc457;
	cam_loc458 <= (internal_wr_en & (internal_wr_ptr == 11'd458) ) ? wr_data : cam_loc458;
	cam_loc459 <= (internal_wr_en & (internal_wr_ptr == 11'd459) ) ? wr_data : cam_loc459;
	cam_loc460 <= (internal_wr_en & (internal_wr_ptr == 11'd460) ) ? wr_data : cam_loc460;
	cam_loc461 <= (internal_wr_en & (internal_wr_ptr == 11'd461) ) ? wr_data : cam_loc461;
	cam_loc462 <= (internal_wr_en & (internal_wr_ptr == 11'd462) ) ? wr_data : cam_loc462;
	cam_loc463 <= (internal_wr_en & (internal_wr_ptr == 11'd463) ) ? wr_data : cam_loc463;
	cam_loc464 <= (internal_wr_en & (internal_wr_ptr == 11'd464) ) ? wr_data : cam_loc464;
	cam_loc465 <= (internal_wr_en & (internal_wr_ptr == 11'd465) ) ? wr_data : cam_loc465;
	cam_loc466 <= (internal_wr_en & (internal_wr_ptr == 11'd466) ) ? wr_data : cam_loc466;
	cam_loc467 <= (internal_wr_en & (internal_wr_ptr == 11'd467) ) ? wr_data : cam_loc467;
	cam_loc468 <= (internal_wr_en & (internal_wr_ptr == 11'd468) ) ? wr_data : cam_loc468;
	cam_loc469 <= (internal_wr_en & (internal_wr_ptr == 11'd469) ) ? wr_data : cam_loc469;
	cam_loc470 <= (internal_wr_en & (internal_wr_ptr == 11'd470) ) ? wr_data : cam_loc470;
	cam_loc471 <= (internal_wr_en & (internal_wr_ptr == 11'd471) ) ? wr_data : cam_loc471;
	cam_loc472 <= (internal_wr_en & (internal_wr_ptr == 11'd472) ) ? wr_data : cam_loc472;
	cam_loc473 <= (internal_wr_en & (internal_wr_ptr == 11'd473) ) ? wr_data : cam_loc473;
	cam_loc474 <= (internal_wr_en & (internal_wr_ptr == 11'd474) ) ? wr_data : cam_loc474;
	cam_loc475 <= (internal_wr_en & (internal_wr_ptr == 11'd475) ) ? wr_data : cam_loc475;
	cam_loc476 <= (internal_wr_en & (internal_wr_ptr == 11'd476) ) ? wr_data : cam_loc476;
	cam_loc477 <= (internal_wr_en & (internal_wr_ptr == 11'd477) ) ? wr_data : cam_loc477;
	cam_loc478 <= (internal_wr_en & (internal_wr_ptr == 11'd478) ) ? wr_data : cam_loc478;
	cam_loc479 <= (internal_wr_en & (internal_wr_ptr == 11'd479) ) ? wr_data : cam_loc479;
	cam_loc480 <= (internal_wr_en & (internal_wr_ptr == 11'd480) ) ? wr_data : cam_loc480;
	cam_loc481 <= (internal_wr_en & (internal_wr_ptr == 11'd481) ) ? wr_data : cam_loc481;
	cam_loc482 <= (internal_wr_en & (internal_wr_ptr == 11'd482) ) ? wr_data : cam_loc482;
	cam_loc483 <= (internal_wr_en & (internal_wr_ptr == 11'd483) ) ? wr_data : cam_loc483;
	cam_loc484 <= (internal_wr_en & (internal_wr_ptr == 11'd484) ) ? wr_data : cam_loc484;
	cam_loc485 <= (internal_wr_en & (internal_wr_ptr == 11'd485) ) ? wr_data : cam_loc485;
	cam_loc486 <= (internal_wr_en & (internal_wr_ptr == 11'd486) ) ? wr_data : cam_loc486;
	cam_loc487 <= (internal_wr_en & (internal_wr_ptr == 11'd487) ) ? wr_data : cam_loc487;
	cam_loc488 <= (internal_wr_en & (internal_wr_ptr == 11'd488) ) ? wr_data : cam_loc488;
	cam_loc489 <= (internal_wr_en & (internal_wr_ptr == 11'd489) ) ? wr_data : cam_loc489;
	cam_loc490 <= (internal_wr_en & (internal_wr_ptr == 11'd490) ) ? wr_data : cam_loc490;
	cam_loc491 <= (internal_wr_en & (internal_wr_ptr == 11'd491) ) ? wr_data : cam_loc491;
	cam_loc492 <= (internal_wr_en & (internal_wr_ptr == 11'd492) ) ? wr_data : cam_loc492;
	cam_loc493 <= (internal_wr_en & (internal_wr_ptr == 11'd493) ) ? wr_data : cam_loc493;
	cam_loc494 <= (internal_wr_en & (internal_wr_ptr == 11'd494) ) ? wr_data : cam_loc494;
	cam_loc495 <= (internal_wr_en & (internal_wr_ptr == 11'd495) ) ? wr_data : cam_loc495;
	cam_loc496 <= (internal_wr_en & (internal_wr_ptr == 11'd496) ) ? wr_data : cam_loc496;
	cam_loc497 <= (internal_wr_en & (internal_wr_ptr == 11'd497) ) ? wr_data : cam_loc497;
	cam_loc498 <= (internal_wr_en & (internal_wr_ptr == 11'd498) ) ? wr_data : cam_loc498;
	cam_loc499 <= (internal_wr_en & (internal_wr_ptr == 11'd499) ) ? wr_data : cam_loc499;
	cam_loc500 <= (internal_wr_en & (internal_wr_ptr == 11'd500) ) ? wr_data : cam_loc500;
	cam_loc501 <= (internal_wr_en & (internal_wr_ptr == 11'd501) ) ? wr_data : cam_loc501;
	cam_loc502 <= (internal_wr_en & (internal_wr_ptr == 11'd502) ) ? wr_data : cam_loc502;
	cam_loc503 <= (internal_wr_en & (internal_wr_ptr == 11'd503) ) ? wr_data : cam_loc503;
	cam_loc504 <= (internal_wr_en & (internal_wr_ptr == 11'd504) ) ? wr_data : cam_loc504;
	cam_loc505 <= (internal_wr_en & (internal_wr_ptr == 11'd505) ) ? wr_data : cam_loc505;
	cam_loc506 <= (internal_wr_en & (internal_wr_ptr == 11'd506) ) ? wr_data : cam_loc506;
	cam_loc507 <= (internal_wr_en & (internal_wr_ptr == 11'd507) ) ? wr_data : cam_loc507;
	cam_loc508 <= (internal_wr_en & (internal_wr_ptr == 11'd508) ) ? wr_data : cam_loc508;
	cam_loc509 <= (internal_wr_en & (internal_wr_ptr == 11'd509) ) ? wr_data : cam_loc509;
	cam_loc510 <= (internal_wr_en & (internal_wr_ptr == 11'd510) ) ? wr_data : cam_loc510;
	cam_loc511 <= (internal_wr_en & (internal_wr_ptr == 11'd511) ) ? wr_data : cam_loc511;
	cam_loc512 <= (internal_wr_en & (internal_wr_ptr == 11'd512) ) ? wr_data : cam_loc512;
	cam_loc513 <= (internal_wr_en & (internal_wr_ptr == 11'd513) ) ? wr_data : cam_loc513;
	cam_loc514 <= (internal_wr_en & (internal_wr_ptr == 11'd514) ) ? wr_data : cam_loc514;
	cam_loc515 <= (internal_wr_en & (internal_wr_ptr == 11'd515) ) ? wr_data : cam_loc515;
	cam_loc516 <= (internal_wr_en & (internal_wr_ptr == 11'd516) ) ? wr_data : cam_loc516;
	cam_loc517 <= (internal_wr_en & (internal_wr_ptr == 11'd517) ) ? wr_data : cam_loc517;
	cam_loc518 <= (internal_wr_en & (internal_wr_ptr == 11'd518) ) ? wr_data : cam_loc518;
	cam_loc519 <= (internal_wr_en & (internal_wr_ptr == 11'd519) ) ? wr_data : cam_loc519;
	cam_loc520 <= (internal_wr_en & (internal_wr_ptr == 11'd520) ) ? wr_data : cam_loc520;
	cam_loc521 <= (internal_wr_en & (internal_wr_ptr == 11'd521) ) ? wr_data : cam_loc521;
	cam_loc522 <= (internal_wr_en & (internal_wr_ptr == 11'd522) ) ? wr_data : cam_loc522;
	cam_loc523 <= (internal_wr_en & (internal_wr_ptr == 11'd523) ) ? wr_data : cam_loc523;
	cam_loc524 <= (internal_wr_en & (internal_wr_ptr == 11'd524) ) ? wr_data : cam_loc524;
	cam_loc525 <= (internal_wr_en & (internal_wr_ptr == 11'd525) ) ? wr_data : cam_loc525;
	cam_loc526 <= (internal_wr_en & (internal_wr_ptr == 11'd526) ) ? wr_data : cam_loc526;
	cam_loc527 <= (internal_wr_en & (internal_wr_ptr == 11'd527) ) ? wr_data : cam_loc527;
	cam_loc528 <= (internal_wr_en & (internal_wr_ptr == 11'd528) ) ? wr_data : cam_loc528;
	cam_loc529 <= (internal_wr_en & (internal_wr_ptr == 11'd529) ) ? wr_data : cam_loc529;
	cam_loc530 <= (internal_wr_en & (internal_wr_ptr == 11'd530) ) ? wr_data : cam_loc530;
	cam_loc531 <= (internal_wr_en & (internal_wr_ptr == 11'd531) ) ? wr_data : cam_loc531;
	cam_loc532 <= (internal_wr_en & (internal_wr_ptr == 11'd532) ) ? wr_data : cam_loc532;
	cam_loc533 <= (internal_wr_en & (internal_wr_ptr == 11'd533) ) ? wr_data : cam_loc533;
	cam_loc534 <= (internal_wr_en & (internal_wr_ptr == 11'd534) ) ? wr_data : cam_loc534;
	cam_loc535 <= (internal_wr_en & (internal_wr_ptr == 11'd535) ) ? wr_data : cam_loc535;
	cam_loc536 <= (internal_wr_en & (internal_wr_ptr == 11'd536) ) ? wr_data : cam_loc536;
	cam_loc537 <= (internal_wr_en & (internal_wr_ptr == 11'd537) ) ? wr_data : cam_loc537;
	cam_loc538 <= (internal_wr_en & (internal_wr_ptr == 11'd538) ) ? wr_data : cam_loc538;
	cam_loc539 <= (internal_wr_en & (internal_wr_ptr == 11'd539) ) ? wr_data : cam_loc539;
	cam_loc540 <= (internal_wr_en & (internal_wr_ptr == 11'd540) ) ? wr_data : cam_loc540;
	cam_loc541 <= (internal_wr_en & (internal_wr_ptr == 11'd541) ) ? wr_data : cam_loc541;
	cam_loc542 <= (internal_wr_en & (internal_wr_ptr == 11'd542) ) ? wr_data : cam_loc542;
	cam_loc543 <= (internal_wr_en & (internal_wr_ptr == 11'd543) ) ? wr_data : cam_loc543;
	cam_loc544 <= (internal_wr_en & (internal_wr_ptr == 11'd544) ) ? wr_data : cam_loc544;
	cam_loc545 <= (internal_wr_en & (internal_wr_ptr == 11'd545) ) ? wr_data : cam_loc545;
	cam_loc546 <= (internal_wr_en & (internal_wr_ptr == 11'd546) ) ? wr_data : cam_loc546;
	cam_loc547 <= (internal_wr_en & (internal_wr_ptr == 11'd547) ) ? wr_data : cam_loc547;
	cam_loc548 <= (internal_wr_en & (internal_wr_ptr == 11'd548) ) ? wr_data : cam_loc548;
	cam_loc549 <= (internal_wr_en & (internal_wr_ptr == 11'd549) ) ? wr_data : cam_loc549;
	cam_loc550 <= (internal_wr_en & (internal_wr_ptr == 11'd550) ) ? wr_data : cam_loc550;
	cam_loc551 <= (internal_wr_en & (internal_wr_ptr == 11'd551) ) ? wr_data : cam_loc551;
	cam_loc552 <= (internal_wr_en & (internal_wr_ptr == 11'd552) ) ? wr_data : cam_loc552;
	cam_loc553 <= (internal_wr_en & (internal_wr_ptr == 11'd553) ) ? wr_data : cam_loc553;
	cam_loc554 <= (internal_wr_en & (internal_wr_ptr == 11'd554) ) ? wr_data : cam_loc554;
	cam_loc555 <= (internal_wr_en & (internal_wr_ptr == 11'd555) ) ? wr_data : cam_loc555;
	cam_loc556 <= (internal_wr_en & (internal_wr_ptr == 11'd556) ) ? wr_data : cam_loc556;
	cam_loc557 <= (internal_wr_en & (internal_wr_ptr == 11'd557) ) ? wr_data : cam_loc557;
	cam_loc558 <= (internal_wr_en & (internal_wr_ptr == 11'd558) ) ? wr_data : cam_loc558;
	cam_loc559 <= (internal_wr_en & (internal_wr_ptr == 11'd559) ) ? wr_data : cam_loc559;
	cam_loc560 <= (internal_wr_en & (internal_wr_ptr == 11'd560) ) ? wr_data : cam_loc560;
	cam_loc561 <= (internal_wr_en & (internal_wr_ptr == 11'd561) ) ? wr_data : cam_loc561;
	cam_loc562 <= (internal_wr_en & (internal_wr_ptr == 11'd562) ) ? wr_data : cam_loc562;
	cam_loc563 <= (internal_wr_en & (internal_wr_ptr == 11'd563) ) ? wr_data : cam_loc563;
	cam_loc564 <= (internal_wr_en & (internal_wr_ptr == 11'd564) ) ? wr_data : cam_loc564;
	cam_loc565 <= (internal_wr_en & (internal_wr_ptr == 11'd565) ) ? wr_data : cam_loc565;
	cam_loc566 <= (internal_wr_en & (internal_wr_ptr == 11'd566) ) ? wr_data : cam_loc566;
	cam_loc567 <= (internal_wr_en & (internal_wr_ptr == 11'd567) ) ? wr_data : cam_loc567;
	cam_loc568 <= (internal_wr_en & (internal_wr_ptr == 11'd568) ) ? wr_data : cam_loc568;
	cam_loc569 <= (internal_wr_en & (internal_wr_ptr == 11'd569) ) ? wr_data : cam_loc569;
	cam_loc570 <= (internal_wr_en & (internal_wr_ptr == 11'd570) ) ? wr_data : cam_loc570;
	cam_loc571 <= (internal_wr_en & (internal_wr_ptr == 11'd571) ) ? wr_data : cam_loc571;
	cam_loc572 <= (internal_wr_en & (internal_wr_ptr == 11'd572) ) ? wr_data : cam_loc572;
	cam_loc573 <= (internal_wr_en & (internal_wr_ptr == 11'd573) ) ? wr_data : cam_loc573;
	cam_loc574 <= (internal_wr_en & (internal_wr_ptr == 11'd574) ) ? wr_data : cam_loc574;
	cam_loc575 <= (internal_wr_en & (internal_wr_ptr == 11'd575) ) ? wr_data : cam_loc575;
	cam_loc576 <= (internal_wr_en & (internal_wr_ptr == 11'd576) ) ? wr_data : cam_loc576;
	cam_loc577 <= (internal_wr_en & (internal_wr_ptr == 11'd577) ) ? wr_data : cam_loc577;
	cam_loc578 <= (internal_wr_en & (internal_wr_ptr == 11'd578) ) ? wr_data : cam_loc578;
	cam_loc579 <= (internal_wr_en & (internal_wr_ptr == 11'd579) ) ? wr_data : cam_loc579;
	cam_loc580 <= (internal_wr_en & (internal_wr_ptr == 11'd580) ) ? wr_data : cam_loc580;
	cam_loc581 <= (internal_wr_en & (internal_wr_ptr == 11'd581) ) ? wr_data : cam_loc581;
	cam_loc582 <= (internal_wr_en & (internal_wr_ptr == 11'd582) ) ? wr_data : cam_loc582;
	cam_loc583 <= (internal_wr_en & (internal_wr_ptr == 11'd583) ) ? wr_data : cam_loc583;
	cam_loc584 <= (internal_wr_en & (internal_wr_ptr == 11'd584) ) ? wr_data : cam_loc584;
	cam_loc585 <= (internal_wr_en & (internal_wr_ptr == 11'd585) ) ? wr_data : cam_loc585;
	cam_loc586 <= (internal_wr_en & (internal_wr_ptr == 11'd586) ) ? wr_data : cam_loc586;
	cam_loc587 <= (internal_wr_en & (internal_wr_ptr == 11'd587) ) ? wr_data : cam_loc587;
	cam_loc588 <= (internal_wr_en & (internal_wr_ptr == 11'd588) ) ? wr_data : cam_loc588;
	cam_loc589 <= (internal_wr_en & (internal_wr_ptr == 11'd589) ) ? wr_data : cam_loc589;
	cam_loc590 <= (internal_wr_en & (internal_wr_ptr == 11'd590) ) ? wr_data : cam_loc590;
	cam_loc591 <= (internal_wr_en & (internal_wr_ptr == 11'd591) ) ? wr_data : cam_loc591;
	cam_loc592 <= (internal_wr_en & (internal_wr_ptr == 11'd592) ) ? wr_data : cam_loc592;
	cam_loc593 <= (internal_wr_en & (internal_wr_ptr == 11'd593) ) ? wr_data : cam_loc593;
	cam_loc594 <= (internal_wr_en & (internal_wr_ptr == 11'd594) ) ? wr_data : cam_loc594;
	cam_loc595 <= (internal_wr_en & (internal_wr_ptr == 11'd595) ) ? wr_data : cam_loc595;
	cam_loc596 <= (internal_wr_en & (internal_wr_ptr == 11'd596) ) ? wr_data : cam_loc596;
	cam_loc597 <= (internal_wr_en & (internal_wr_ptr == 11'd597) ) ? wr_data : cam_loc597;
	cam_loc598 <= (internal_wr_en & (internal_wr_ptr == 11'd598) ) ? wr_data : cam_loc598;
	cam_loc599 <= (internal_wr_en & (internal_wr_ptr == 11'd599) ) ? wr_data : cam_loc599;
	cam_loc600 <= (internal_wr_en & (internal_wr_ptr == 11'd600) ) ? wr_data : cam_loc600;
	cam_loc601 <= (internal_wr_en & (internal_wr_ptr == 11'd601) ) ? wr_data : cam_loc601;
	cam_loc602 <= (internal_wr_en & (internal_wr_ptr == 11'd602) ) ? wr_data : cam_loc602;
	cam_loc603 <= (internal_wr_en & (internal_wr_ptr == 11'd603) ) ? wr_data : cam_loc603;
	cam_loc604 <= (internal_wr_en & (internal_wr_ptr == 11'd604) ) ? wr_data : cam_loc604;
	cam_loc605 <= (internal_wr_en & (internal_wr_ptr == 11'd605) ) ? wr_data : cam_loc605;
	cam_loc606 <= (internal_wr_en & (internal_wr_ptr == 11'd606) ) ? wr_data : cam_loc606;
	cam_loc607 <= (internal_wr_en & (internal_wr_ptr == 11'd607) ) ? wr_data : cam_loc607;
	cam_loc608 <= (internal_wr_en & (internal_wr_ptr == 11'd608) ) ? wr_data : cam_loc608;
	cam_loc609 <= (internal_wr_en & (internal_wr_ptr == 11'd609) ) ? wr_data : cam_loc609;
	cam_loc610 <= (internal_wr_en & (internal_wr_ptr == 11'd610) ) ? wr_data : cam_loc610;
	cam_loc611 <= (internal_wr_en & (internal_wr_ptr == 11'd611) ) ? wr_data : cam_loc611;
	cam_loc612 <= (internal_wr_en & (internal_wr_ptr == 11'd612) ) ? wr_data : cam_loc612;
	cam_loc613 <= (internal_wr_en & (internal_wr_ptr == 11'd613) ) ? wr_data : cam_loc613;
	cam_loc614 <= (internal_wr_en & (internal_wr_ptr == 11'd614) ) ? wr_data : cam_loc614;
	cam_loc615 <= (internal_wr_en & (internal_wr_ptr == 11'd615) ) ? wr_data : cam_loc615;
	cam_loc616 <= (internal_wr_en & (internal_wr_ptr == 11'd616) ) ? wr_data : cam_loc616;
	cam_loc617 <= (internal_wr_en & (internal_wr_ptr == 11'd617) ) ? wr_data : cam_loc617;
	cam_loc618 <= (internal_wr_en & (internal_wr_ptr == 11'd618) ) ? wr_data : cam_loc618;
	cam_loc619 <= (internal_wr_en & (internal_wr_ptr == 11'd619) ) ? wr_data : cam_loc619;
	cam_loc620 <= (internal_wr_en & (internal_wr_ptr == 11'd620) ) ? wr_data : cam_loc620;
	cam_loc621 <= (internal_wr_en & (internal_wr_ptr == 11'd621) ) ? wr_data : cam_loc621;
	cam_loc622 <= (internal_wr_en & (internal_wr_ptr == 11'd622) ) ? wr_data : cam_loc622;
	cam_loc623 <= (internal_wr_en & (internal_wr_ptr == 11'd623) ) ? wr_data : cam_loc623;
	cam_loc624 <= (internal_wr_en & (internal_wr_ptr == 11'd624) ) ? wr_data : cam_loc624;
	cam_loc625 <= (internal_wr_en & (internal_wr_ptr == 11'd625) ) ? wr_data : cam_loc625;
	cam_loc626 <= (internal_wr_en & (internal_wr_ptr == 11'd626) ) ? wr_data : cam_loc626;
	cam_loc627 <= (internal_wr_en & (internal_wr_ptr == 11'd627) ) ? wr_data : cam_loc627;
	cam_loc628 <= (internal_wr_en & (internal_wr_ptr == 11'd628) ) ? wr_data : cam_loc628;
	cam_loc629 <= (internal_wr_en & (internal_wr_ptr == 11'd629) ) ? wr_data : cam_loc629;
	cam_loc630 <= (internal_wr_en & (internal_wr_ptr == 11'd630) ) ? wr_data : cam_loc630;
	cam_loc631 <= (internal_wr_en & (internal_wr_ptr == 11'd631) ) ? wr_data : cam_loc631;
	cam_loc632 <= (internal_wr_en & (internal_wr_ptr == 11'd632) ) ? wr_data : cam_loc632;
	cam_loc633 <= (internal_wr_en & (internal_wr_ptr == 11'd633) ) ? wr_data : cam_loc633;
	cam_loc634 <= (internal_wr_en & (internal_wr_ptr == 11'd634) ) ? wr_data : cam_loc634;
	cam_loc635 <= (internal_wr_en & (internal_wr_ptr == 11'd635) ) ? wr_data : cam_loc635;
	cam_loc636 <= (internal_wr_en & (internal_wr_ptr == 11'd636) ) ? wr_data : cam_loc636;
	cam_loc637 <= (internal_wr_en & (internal_wr_ptr == 11'd637) ) ? wr_data : cam_loc637;
	cam_loc638 <= (internal_wr_en & (internal_wr_ptr == 11'd638) ) ? wr_data : cam_loc638;
	cam_loc639 <= (internal_wr_en & (internal_wr_ptr == 11'd639) ) ? wr_data : cam_loc639;
	cam_loc640 <= (internal_wr_en & (internal_wr_ptr == 11'd640) ) ? wr_data : cam_loc640;
	cam_loc641 <= (internal_wr_en & (internal_wr_ptr == 11'd641) ) ? wr_data : cam_loc641;
	cam_loc642 <= (internal_wr_en & (internal_wr_ptr == 11'd642) ) ? wr_data : cam_loc642;
	cam_loc643 <= (internal_wr_en & (internal_wr_ptr == 11'd643) ) ? wr_data : cam_loc643;
	cam_loc644 <= (internal_wr_en & (internal_wr_ptr == 11'd644) ) ? wr_data : cam_loc644;
	cam_loc645 <= (internal_wr_en & (internal_wr_ptr == 11'd645) ) ? wr_data : cam_loc645;
	cam_loc646 <= (internal_wr_en & (internal_wr_ptr == 11'd646) ) ? wr_data : cam_loc646;
	cam_loc647 <= (internal_wr_en & (internal_wr_ptr == 11'd647) ) ? wr_data : cam_loc647;
	cam_loc648 <= (internal_wr_en & (internal_wr_ptr == 11'd648) ) ? wr_data : cam_loc648;
	cam_loc649 <= (internal_wr_en & (internal_wr_ptr == 11'd649) ) ? wr_data : cam_loc649;
	cam_loc650 <= (internal_wr_en & (internal_wr_ptr == 11'd650) ) ? wr_data : cam_loc650;
	cam_loc651 <= (internal_wr_en & (internal_wr_ptr == 11'd651) ) ? wr_data : cam_loc651;
	cam_loc652 <= (internal_wr_en & (internal_wr_ptr == 11'd652) ) ? wr_data : cam_loc652;
	cam_loc653 <= (internal_wr_en & (internal_wr_ptr == 11'd653) ) ? wr_data : cam_loc653;
	cam_loc654 <= (internal_wr_en & (internal_wr_ptr == 11'd654) ) ? wr_data : cam_loc654;
	cam_loc655 <= (internal_wr_en & (internal_wr_ptr == 11'd655) ) ? wr_data : cam_loc655;
	cam_loc656 <= (internal_wr_en & (internal_wr_ptr == 11'd656) ) ? wr_data : cam_loc656;
	cam_loc657 <= (internal_wr_en & (internal_wr_ptr == 11'd657) ) ? wr_data : cam_loc657;
	cam_loc658 <= (internal_wr_en & (internal_wr_ptr == 11'd658) ) ? wr_data : cam_loc658;
	cam_loc659 <= (internal_wr_en & (internal_wr_ptr == 11'd659) ) ? wr_data : cam_loc659;
	cam_loc660 <= (internal_wr_en & (internal_wr_ptr == 11'd660) ) ? wr_data : cam_loc660;
	cam_loc661 <= (internal_wr_en & (internal_wr_ptr == 11'd661) ) ? wr_data : cam_loc661;
	cam_loc662 <= (internal_wr_en & (internal_wr_ptr == 11'd662) ) ? wr_data : cam_loc662;
	cam_loc663 <= (internal_wr_en & (internal_wr_ptr == 11'd663) ) ? wr_data : cam_loc663;
	cam_loc664 <= (internal_wr_en & (internal_wr_ptr == 11'd664) ) ? wr_data : cam_loc664;
	cam_loc665 <= (internal_wr_en & (internal_wr_ptr == 11'd665) ) ? wr_data : cam_loc665;
	cam_loc666 <= (internal_wr_en & (internal_wr_ptr == 11'd666) ) ? wr_data : cam_loc666;
	cam_loc667 <= (internal_wr_en & (internal_wr_ptr == 11'd667) ) ? wr_data : cam_loc667;
	cam_loc668 <= (internal_wr_en & (internal_wr_ptr == 11'd668) ) ? wr_data : cam_loc668;
	cam_loc669 <= (internal_wr_en & (internal_wr_ptr == 11'd669) ) ? wr_data : cam_loc669;
	cam_loc670 <= (internal_wr_en & (internal_wr_ptr == 11'd670) ) ? wr_data : cam_loc670;
	cam_loc671 <= (internal_wr_en & (internal_wr_ptr == 11'd671) ) ? wr_data : cam_loc671;
	cam_loc672 <= (internal_wr_en & (internal_wr_ptr == 11'd672) ) ? wr_data : cam_loc672;
	cam_loc673 <= (internal_wr_en & (internal_wr_ptr == 11'd673) ) ? wr_data : cam_loc673;
	cam_loc674 <= (internal_wr_en & (internal_wr_ptr == 11'd674) ) ? wr_data : cam_loc674;
	cam_loc675 <= (internal_wr_en & (internal_wr_ptr == 11'd675) ) ? wr_data : cam_loc675;
	cam_loc676 <= (internal_wr_en & (internal_wr_ptr == 11'd676) ) ? wr_data : cam_loc676;
	cam_loc677 <= (internal_wr_en & (internal_wr_ptr == 11'd677) ) ? wr_data : cam_loc677;
	cam_loc678 <= (internal_wr_en & (internal_wr_ptr == 11'd678) ) ? wr_data : cam_loc678;
	cam_loc679 <= (internal_wr_en & (internal_wr_ptr == 11'd679) ) ? wr_data : cam_loc679;
	cam_loc680 <= (internal_wr_en & (internal_wr_ptr == 11'd680) ) ? wr_data : cam_loc680;
	cam_loc681 <= (internal_wr_en & (internal_wr_ptr == 11'd681) ) ? wr_data : cam_loc681;
	cam_loc682 <= (internal_wr_en & (internal_wr_ptr == 11'd682) ) ? wr_data : cam_loc682;
	cam_loc683 <= (internal_wr_en & (internal_wr_ptr == 11'd683) ) ? wr_data : cam_loc683;
	cam_loc684 <= (internal_wr_en & (internal_wr_ptr == 11'd684) ) ? wr_data : cam_loc684;
	cam_loc685 <= (internal_wr_en & (internal_wr_ptr == 11'd685) ) ? wr_data : cam_loc685;
	cam_loc686 <= (internal_wr_en & (internal_wr_ptr == 11'd686) ) ? wr_data : cam_loc686;
	cam_loc687 <= (internal_wr_en & (internal_wr_ptr == 11'd687) ) ? wr_data : cam_loc687;
	cam_loc688 <= (internal_wr_en & (internal_wr_ptr == 11'd688) ) ? wr_data : cam_loc688;
	cam_loc689 <= (internal_wr_en & (internal_wr_ptr == 11'd689) ) ? wr_data : cam_loc689;
	cam_loc690 <= (internal_wr_en & (internal_wr_ptr == 11'd690) ) ? wr_data : cam_loc690;
	cam_loc691 <= (internal_wr_en & (internal_wr_ptr == 11'd691) ) ? wr_data : cam_loc691;
	cam_loc692 <= (internal_wr_en & (internal_wr_ptr == 11'd692) ) ? wr_data : cam_loc692;
	cam_loc693 <= (internal_wr_en & (internal_wr_ptr == 11'd693) ) ? wr_data : cam_loc693;
	cam_loc694 <= (internal_wr_en & (internal_wr_ptr == 11'd694) ) ? wr_data : cam_loc694;
	cam_loc695 <= (internal_wr_en & (internal_wr_ptr == 11'd695) ) ? wr_data : cam_loc695;
	cam_loc696 <= (internal_wr_en & (internal_wr_ptr == 11'd696) ) ? wr_data : cam_loc696;
	cam_loc697 <= (internal_wr_en & (internal_wr_ptr == 11'd697) ) ? wr_data : cam_loc697;
	cam_loc698 <= (internal_wr_en & (internal_wr_ptr == 11'd698) ) ? wr_data : cam_loc698;
	cam_loc699 <= (internal_wr_en & (internal_wr_ptr == 11'd699) ) ? wr_data : cam_loc699;
	cam_loc700 <= (internal_wr_en & (internal_wr_ptr == 11'd700) ) ? wr_data : cam_loc700;
	cam_loc701 <= (internal_wr_en & (internal_wr_ptr == 11'd701) ) ? wr_data : cam_loc701;
	cam_loc702 <= (internal_wr_en & (internal_wr_ptr == 11'd702) ) ? wr_data : cam_loc702;
	cam_loc703 <= (internal_wr_en & (internal_wr_ptr == 11'd703) ) ? wr_data : cam_loc703;
	cam_loc704 <= (internal_wr_en & (internal_wr_ptr == 11'd704) ) ? wr_data : cam_loc704;
	cam_loc705 <= (internal_wr_en & (internal_wr_ptr == 11'd705) ) ? wr_data : cam_loc705;
	cam_loc706 <= (internal_wr_en & (internal_wr_ptr == 11'd706) ) ? wr_data : cam_loc706;
	cam_loc707 <= (internal_wr_en & (internal_wr_ptr == 11'd707) ) ? wr_data : cam_loc707;
	cam_loc708 <= (internal_wr_en & (internal_wr_ptr == 11'd708) ) ? wr_data : cam_loc708;
	cam_loc709 <= (internal_wr_en & (internal_wr_ptr == 11'd709) ) ? wr_data : cam_loc709;
	cam_loc710 <= (internal_wr_en & (internal_wr_ptr == 11'd710) ) ? wr_data : cam_loc710;
	cam_loc711 <= (internal_wr_en & (internal_wr_ptr == 11'd711) ) ? wr_data : cam_loc711;
	cam_loc712 <= (internal_wr_en & (internal_wr_ptr == 11'd712) ) ? wr_data : cam_loc712;
	cam_loc713 <= (internal_wr_en & (internal_wr_ptr == 11'd713) ) ? wr_data : cam_loc713;
	cam_loc714 <= (internal_wr_en & (internal_wr_ptr == 11'd714) ) ? wr_data : cam_loc714;
	cam_loc715 <= (internal_wr_en & (internal_wr_ptr == 11'd715) ) ? wr_data : cam_loc715;
	cam_loc716 <= (internal_wr_en & (internal_wr_ptr == 11'd716) ) ? wr_data : cam_loc716;
	cam_loc717 <= (internal_wr_en & (internal_wr_ptr == 11'd717) ) ? wr_data : cam_loc717;
	cam_loc718 <= (internal_wr_en & (internal_wr_ptr == 11'd718) ) ? wr_data : cam_loc718;
	cam_loc719 <= (internal_wr_en & (internal_wr_ptr == 11'd719) ) ? wr_data : cam_loc719;
	cam_loc720 <= (internal_wr_en & (internal_wr_ptr == 11'd720) ) ? wr_data : cam_loc720;
	cam_loc721 <= (internal_wr_en & (internal_wr_ptr == 11'd721) ) ? wr_data : cam_loc721;
	cam_loc722 <= (internal_wr_en & (internal_wr_ptr == 11'd722) ) ? wr_data : cam_loc722;
	cam_loc723 <= (internal_wr_en & (internal_wr_ptr == 11'd723) ) ? wr_data : cam_loc723;
	cam_loc724 <= (internal_wr_en & (internal_wr_ptr == 11'd724) ) ? wr_data : cam_loc724;
	cam_loc725 <= (internal_wr_en & (internal_wr_ptr == 11'd725) ) ? wr_data : cam_loc725;
	cam_loc726 <= (internal_wr_en & (internal_wr_ptr == 11'd726) ) ? wr_data : cam_loc726;
	cam_loc727 <= (internal_wr_en & (internal_wr_ptr == 11'd727) ) ? wr_data : cam_loc727;
	cam_loc728 <= (internal_wr_en & (internal_wr_ptr == 11'd728) ) ? wr_data : cam_loc728;
	cam_loc729 <= (internal_wr_en & (internal_wr_ptr == 11'd729) ) ? wr_data : cam_loc729;
	cam_loc730 <= (internal_wr_en & (internal_wr_ptr == 11'd730) ) ? wr_data : cam_loc730;
	cam_loc731 <= (internal_wr_en & (internal_wr_ptr == 11'd731) ) ? wr_data : cam_loc731;
	cam_loc732 <= (internal_wr_en & (internal_wr_ptr == 11'd732) ) ? wr_data : cam_loc732;
	cam_loc733 <= (internal_wr_en & (internal_wr_ptr == 11'd733) ) ? wr_data : cam_loc733;
	cam_loc734 <= (internal_wr_en & (internal_wr_ptr == 11'd734) ) ? wr_data : cam_loc734;
	cam_loc735 <= (internal_wr_en & (internal_wr_ptr == 11'd735) ) ? wr_data : cam_loc735;
	cam_loc736 <= (internal_wr_en & (internal_wr_ptr == 11'd736) ) ? wr_data : cam_loc736;
	cam_loc737 <= (internal_wr_en & (internal_wr_ptr == 11'd737) ) ? wr_data : cam_loc737;
	cam_loc738 <= (internal_wr_en & (internal_wr_ptr == 11'd738) ) ? wr_data : cam_loc738;
	cam_loc739 <= (internal_wr_en & (internal_wr_ptr == 11'd739) ) ? wr_data : cam_loc739;
	cam_loc740 <= (internal_wr_en & (internal_wr_ptr == 11'd740) ) ? wr_data : cam_loc740;
	cam_loc741 <= (internal_wr_en & (internal_wr_ptr == 11'd741) ) ? wr_data : cam_loc741;
	cam_loc742 <= (internal_wr_en & (internal_wr_ptr == 11'd742) ) ? wr_data : cam_loc742;
	cam_loc743 <= (internal_wr_en & (internal_wr_ptr == 11'd743) ) ? wr_data : cam_loc743;
	cam_loc744 <= (internal_wr_en & (internal_wr_ptr == 11'd744) ) ? wr_data : cam_loc744;
	cam_loc745 <= (internal_wr_en & (internal_wr_ptr == 11'd745) ) ? wr_data : cam_loc745;
	cam_loc746 <= (internal_wr_en & (internal_wr_ptr == 11'd746) ) ? wr_data : cam_loc746;
	cam_loc747 <= (internal_wr_en & (internal_wr_ptr == 11'd747) ) ? wr_data : cam_loc747;
	cam_loc748 <= (internal_wr_en & (internal_wr_ptr == 11'd748) ) ? wr_data : cam_loc748;
	cam_loc749 <= (internal_wr_en & (internal_wr_ptr == 11'd749) ) ? wr_data : cam_loc749;
	cam_loc750 <= (internal_wr_en & (internal_wr_ptr == 11'd750) ) ? wr_data : cam_loc750;
	cam_loc751 <= (internal_wr_en & (internal_wr_ptr == 11'd751) ) ? wr_data : cam_loc751;
	cam_loc752 <= (internal_wr_en & (internal_wr_ptr == 11'd752) ) ? wr_data : cam_loc752;
	cam_loc753 <= (internal_wr_en & (internal_wr_ptr == 11'd753) ) ? wr_data : cam_loc753;
	cam_loc754 <= (internal_wr_en & (internal_wr_ptr == 11'd754) ) ? wr_data : cam_loc754;
	cam_loc755 <= (internal_wr_en & (internal_wr_ptr == 11'd755) ) ? wr_data : cam_loc755;
	cam_loc756 <= (internal_wr_en & (internal_wr_ptr == 11'd756) ) ? wr_data : cam_loc756;
	cam_loc757 <= (internal_wr_en & (internal_wr_ptr == 11'd757) ) ? wr_data : cam_loc757;
	cam_loc758 <= (internal_wr_en & (internal_wr_ptr == 11'd758) ) ? wr_data : cam_loc758;
	cam_loc759 <= (internal_wr_en & (internal_wr_ptr == 11'd759) ) ? wr_data : cam_loc759;
	cam_loc760 <= (internal_wr_en & (internal_wr_ptr == 11'd760) ) ? wr_data : cam_loc760;
	cam_loc761 <= (internal_wr_en & (internal_wr_ptr == 11'd761) ) ? wr_data : cam_loc761;
	cam_loc762 <= (internal_wr_en & (internal_wr_ptr == 11'd762) ) ? wr_data : cam_loc762;
	cam_loc763 <= (internal_wr_en & (internal_wr_ptr == 11'd763) ) ? wr_data : cam_loc763;
	cam_loc764 <= (internal_wr_en & (internal_wr_ptr == 11'd764) ) ? wr_data : cam_loc764;
	cam_loc765 <= (internal_wr_en & (internal_wr_ptr == 11'd765) ) ? wr_data : cam_loc765;
	cam_loc766 <= (internal_wr_en & (internal_wr_ptr == 11'd766) ) ? wr_data : cam_loc766;
	cam_loc767 <= (internal_wr_en & (internal_wr_ptr == 11'd767) ) ? wr_data : cam_loc767;
	cam_loc768 <= (internal_wr_en & (internal_wr_ptr == 11'd768) ) ? wr_data : cam_loc768;
	cam_loc769 <= (internal_wr_en & (internal_wr_ptr == 11'd769) ) ? wr_data : cam_loc769;
	cam_loc770 <= (internal_wr_en & (internal_wr_ptr == 11'd770) ) ? wr_data : cam_loc770;
	cam_loc771 <= (internal_wr_en & (internal_wr_ptr == 11'd771) ) ? wr_data : cam_loc771;
	cam_loc772 <= (internal_wr_en & (internal_wr_ptr == 11'd772) ) ? wr_data : cam_loc772;
	cam_loc773 <= (internal_wr_en & (internal_wr_ptr == 11'd773) ) ? wr_data : cam_loc773;
	cam_loc774 <= (internal_wr_en & (internal_wr_ptr == 11'd774) ) ? wr_data : cam_loc774;
	cam_loc775 <= (internal_wr_en & (internal_wr_ptr == 11'd775) ) ? wr_data : cam_loc775;
	cam_loc776 <= (internal_wr_en & (internal_wr_ptr == 11'd776) ) ? wr_data : cam_loc776;
	cam_loc777 <= (internal_wr_en & (internal_wr_ptr == 11'd777) ) ? wr_data : cam_loc777;
	cam_loc778 <= (internal_wr_en & (internal_wr_ptr == 11'd778) ) ? wr_data : cam_loc778;
	cam_loc779 <= (internal_wr_en & (internal_wr_ptr == 11'd779) ) ? wr_data : cam_loc779;
	cam_loc780 <= (internal_wr_en & (internal_wr_ptr == 11'd780) ) ? wr_data : cam_loc780;
	cam_loc781 <= (internal_wr_en & (internal_wr_ptr == 11'd781) ) ? wr_data : cam_loc781;
	cam_loc782 <= (internal_wr_en & (internal_wr_ptr == 11'd782) ) ? wr_data : cam_loc782;
	cam_loc783 <= (internal_wr_en & (internal_wr_ptr == 11'd783) ) ? wr_data : cam_loc783;
	cam_loc784 <= (internal_wr_en & (internal_wr_ptr == 11'd784) ) ? wr_data : cam_loc784;
	cam_loc785 <= (internal_wr_en & (internal_wr_ptr == 11'd785) ) ? wr_data : cam_loc785;
	cam_loc786 <= (internal_wr_en & (internal_wr_ptr == 11'd786) ) ? wr_data : cam_loc786;
	cam_loc787 <= (internal_wr_en & (internal_wr_ptr == 11'd787) ) ? wr_data : cam_loc787;
	cam_loc788 <= (internal_wr_en & (internal_wr_ptr == 11'd788) ) ? wr_data : cam_loc788;
	cam_loc789 <= (internal_wr_en & (internal_wr_ptr == 11'd789) ) ? wr_data : cam_loc789;
	cam_loc790 <= (internal_wr_en & (internal_wr_ptr == 11'd790) ) ? wr_data : cam_loc790;
	cam_loc791 <= (internal_wr_en & (internal_wr_ptr == 11'd791) ) ? wr_data : cam_loc791;
	cam_loc792 <= (internal_wr_en & (internal_wr_ptr == 11'd792) ) ? wr_data : cam_loc792;
	cam_loc793 <= (internal_wr_en & (internal_wr_ptr == 11'd793) ) ? wr_data : cam_loc793;
	cam_loc794 <= (internal_wr_en & (internal_wr_ptr == 11'd794) ) ? wr_data : cam_loc794;
	cam_loc795 <= (internal_wr_en & (internal_wr_ptr == 11'd795) ) ? wr_data : cam_loc795;
	cam_loc796 <= (internal_wr_en & (internal_wr_ptr == 11'd796) ) ? wr_data : cam_loc796;
	cam_loc797 <= (internal_wr_en & (internal_wr_ptr == 11'd797) ) ? wr_data : cam_loc797;
	cam_loc798 <= (internal_wr_en & (internal_wr_ptr == 11'd798) ) ? wr_data : cam_loc798;
	cam_loc799 <= (internal_wr_en & (internal_wr_ptr == 11'd799) ) ? wr_data : cam_loc799;
	cam_loc800 <= (internal_wr_en & (internal_wr_ptr == 11'd800) ) ? wr_data : cam_loc800;
	cam_loc801 <= (internal_wr_en & (internal_wr_ptr == 11'd801) ) ? wr_data : cam_loc801;
	cam_loc802 <= (internal_wr_en & (internal_wr_ptr == 11'd802) ) ? wr_data : cam_loc802;
	cam_loc803 <= (internal_wr_en & (internal_wr_ptr == 11'd803) ) ? wr_data : cam_loc803;
	cam_loc804 <= (internal_wr_en & (internal_wr_ptr == 11'd804) ) ? wr_data : cam_loc804;
	cam_loc805 <= (internal_wr_en & (internal_wr_ptr == 11'd805) ) ? wr_data : cam_loc805;
	cam_loc806 <= (internal_wr_en & (internal_wr_ptr == 11'd806) ) ? wr_data : cam_loc806;
	cam_loc807 <= (internal_wr_en & (internal_wr_ptr == 11'd807) ) ? wr_data : cam_loc807;
	cam_loc808 <= (internal_wr_en & (internal_wr_ptr == 11'd808) ) ? wr_data : cam_loc808;
	cam_loc809 <= (internal_wr_en & (internal_wr_ptr == 11'd809) ) ? wr_data : cam_loc809;
	cam_loc810 <= (internal_wr_en & (internal_wr_ptr == 11'd810) ) ? wr_data : cam_loc810;
	cam_loc811 <= (internal_wr_en & (internal_wr_ptr == 11'd811) ) ? wr_data : cam_loc811;
	cam_loc812 <= (internal_wr_en & (internal_wr_ptr == 11'd812) ) ? wr_data : cam_loc812;
	cam_loc813 <= (internal_wr_en & (internal_wr_ptr == 11'd813) ) ? wr_data : cam_loc813;
	cam_loc814 <= (internal_wr_en & (internal_wr_ptr == 11'd814) ) ? wr_data : cam_loc814;
	cam_loc815 <= (internal_wr_en & (internal_wr_ptr == 11'd815) ) ? wr_data : cam_loc815;
	cam_loc816 <= (internal_wr_en & (internal_wr_ptr == 11'd816) ) ? wr_data : cam_loc816;
	cam_loc817 <= (internal_wr_en & (internal_wr_ptr == 11'd817) ) ? wr_data : cam_loc817;
	cam_loc818 <= (internal_wr_en & (internal_wr_ptr == 11'd818) ) ? wr_data : cam_loc818;
	cam_loc819 <= (internal_wr_en & (internal_wr_ptr == 11'd819) ) ? wr_data : cam_loc819;
	cam_loc820 <= (internal_wr_en & (internal_wr_ptr == 11'd820) ) ? wr_data : cam_loc820;
	cam_loc821 <= (internal_wr_en & (internal_wr_ptr == 11'd821) ) ? wr_data : cam_loc821;
	cam_loc822 <= (internal_wr_en & (internal_wr_ptr == 11'd822) ) ? wr_data : cam_loc822;
	cam_loc823 <= (internal_wr_en & (internal_wr_ptr == 11'd823) ) ? wr_data : cam_loc823;
	cam_loc824 <= (internal_wr_en & (internal_wr_ptr == 11'd824) ) ? wr_data : cam_loc824;
	cam_loc825 <= (internal_wr_en & (internal_wr_ptr == 11'd825) ) ? wr_data : cam_loc825;
	cam_loc826 <= (internal_wr_en & (internal_wr_ptr == 11'd826) ) ? wr_data : cam_loc826;
	cam_loc827 <= (internal_wr_en & (internal_wr_ptr == 11'd827) ) ? wr_data : cam_loc827;
	cam_loc828 <= (internal_wr_en & (internal_wr_ptr == 11'd828) ) ? wr_data : cam_loc828;
	cam_loc829 <= (internal_wr_en & (internal_wr_ptr == 11'd829) ) ? wr_data : cam_loc829;
	cam_loc830 <= (internal_wr_en & (internal_wr_ptr == 11'd830) ) ? wr_data : cam_loc830;
	cam_loc831 <= (internal_wr_en & (internal_wr_ptr == 11'd831) ) ? wr_data : cam_loc831;
	cam_loc832 <= (internal_wr_en & (internal_wr_ptr == 11'd832) ) ? wr_data : cam_loc832;
	cam_loc833 <= (internal_wr_en & (internal_wr_ptr == 11'd833) ) ? wr_data : cam_loc833;
	cam_loc834 <= (internal_wr_en & (internal_wr_ptr == 11'd834) ) ? wr_data : cam_loc834;
	cam_loc835 <= (internal_wr_en & (internal_wr_ptr == 11'd835) ) ? wr_data : cam_loc835;
	cam_loc836 <= (internal_wr_en & (internal_wr_ptr == 11'd836) ) ? wr_data : cam_loc836;
	cam_loc837 <= (internal_wr_en & (internal_wr_ptr == 11'd837) ) ? wr_data : cam_loc837;
	cam_loc838 <= (internal_wr_en & (internal_wr_ptr == 11'd838) ) ? wr_data : cam_loc838;
	cam_loc839 <= (internal_wr_en & (internal_wr_ptr == 11'd839) ) ? wr_data : cam_loc839;
	cam_loc840 <= (internal_wr_en & (internal_wr_ptr == 11'd840) ) ? wr_data : cam_loc840;
	cam_loc841 <= (internal_wr_en & (internal_wr_ptr == 11'd841) ) ? wr_data : cam_loc841;
	cam_loc842 <= (internal_wr_en & (internal_wr_ptr == 11'd842) ) ? wr_data : cam_loc842;
	cam_loc843 <= (internal_wr_en & (internal_wr_ptr == 11'd843) ) ? wr_data : cam_loc843;
	cam_loc844 <= (internal_wr_en & (internal_wr_ptr == 11'd844) ) ? wr_data : cam_loc844;
	cam_loc845 <= (internal_wr_en & (internal_wr_ptr == 11'd845) ) ? wr_data : cam_loc845;
	cam_loc846 <= (internal_wr_en & (internal_wr_ptr == 11'd846) ) ? wr_data : cam_loc846;
	cam_loc847 <= (internal_wr_en & (internal_wr_ptr == 11'd847) ) ? wr_data : cam_loc847;
	cam_loc848 <= (internal_wr_en & (internal_wr_ptr == 11'd848) ) ? wr_data : cam_loc848;
	cam_loc849 <= (internal_wr_en & (internal_wr_ptr == 11'd849) ) ? wr_data : cam_loc849;
	cam_loc850 <= (internal_wr_en & (internal_wr_ptr == 11'd850) ) ? wr_data : cam_loc850;
	cam_loc851 <= (internal_wr_en & (internal_wr_ptr == 11'd851) ) ? wr_data : cam_loc851;
	cam_loc852 <= (internal_wr_en & (internal_wr_ptr == 11'd852) ) ? wr_data : cam_loc852;
	cam_loc853 <= (internal_wr_en & (internal_wr_ptr == 11'd853) ) ? wr_data : cam_loc853;
	cam_loc854 <= (internal_wr_en & (internal_wr_ptr == 11'd854) ) ? wr_data : cam_loc854;
	cam_loc855 <= (internal_wr_en & (internal_wr_ptr == 11'd855) ) ? wr_data : cam_loc855;
	cam_loc856 <= (internal_wr_en & (internal_wr_ptr == 11'd856) ) ? wr_data : cam_loc856;
	cam_loc857 <= (internal_wr_en & (internal_wr_ptr == 11'd857) ) ? wr_data : cam_loc857;
	cam_loc858 <= (internal_wr_en & (internal_wr_ptr == 11'd858) ) ? wr_data : cam_loc858;
	cam_loc859 <= (internal_wr_en & (internal_wr_ptr == 11'd859) ) ? wr_data : cam_loc859;
	cam_loc860 <= (internal_wr_en & (internal_wr_ptr == 11'd860) ) ? wr_data : cam_loc860;
	cam_loc861 <= (internal_wr_en & (internal_wr_ptr == 11'd861) ) ? wr_data : cam_loc861;
	cam_loc862 <= (internal_wr_en & (internal_wr_ptr == 11'd862) ) ? wr_data : cam_loc862;
	cam_loc863 <= (internal_wr_en & (internal_wr_ptr == 11'd863) ) ? wr_data : cam_loc863;
	cam_loc864 <= (internal_wr_en & (internal_wr_ptr == 11'd864) ) ? wr_data : cam_loc864;
	cam_loc865 <= (internal_wr_en & (internal_wr_ptr == 11'd865) ) ? wr_data : cam_loc865;
	cam_loc866 <= (internal_wr_en & (internal_wr_ptr == 11'd866) ) ? wr_data : cam_loc866;
	cam_loc867 <= (internal_wr_en & (internal_wr_ptr == 11'd867) ) ? wr_data : cam_loc867;
	cam_loc868 <= (internal_wr_en & (internal_wr_ptr == 11'd868) ) ? wr_data : cam_loc868;
	cam_loc869 <= (internal_wr_en & (internal_wr_ptr == 11'd869) ) ? wr_data : cam_loc869;
	cam_loc870 <= (internal_wr_en & (internal_wr_ptr == 11'd870) ) ? wr_data : cam_loc870;
	cam_loc871 <= (internal_wr_en & (internal_wr_ptr == 11'd871) ) ? wr_data : cam_loc871;
	cam_loc872 <= (internal_wr_en & (internal_wr_ptr == 11'd872) ) ? wr_data : cam_loc872;
	cam_loc873 <= (internal_wr_en & (internal_wr_ptr == 11'd873) ) ? wr_data : cam_loc873;
	cam_loc874 <= (internal_wr_en & (internal_wr_ptr == 11'd874) ) ? wr_data : cam_loc874;
	cam_loc875 <= (internal_wr_en & (internal_wr_ptr == 11'd875) ) ? wr_data : cam_loc875;
	cam_loc876 <= (internal_wr_en & (internal_wr_ptr == 11'd876) ) ? wr_data : cam_loc876;
	cam_loc877 <= (internal_wr_en & (internal_wr_ptr == 11'd877) ) ? wr_data : cam_loc877;
	cam_loc878 <= (internal_wr_en & (internal_wr_ptr == 11'd878) ) ? wr_data : cam_loc878;
	cam_loc879 <= (internal_wr_en & (internal_wr_ptr == 11'd879) ) ? wr_data : cam_loc879;
	cam_loc880 <= (internal_wr_en & (internal_wr_ptr == 11'd880) ) ? wr_data : cam_loc880;
	cam_loc881 <= (internal_wr_en & (internal_wr_ptr == 11'd881) ) ? wr_data : cam_loc881;
	cam_loc882 <= (internal_wr_en & (internal_wr_ptr == 11'd882) ) ? wr_data : cam_loc882;
	cam_loc883 <= (internal_wr_en & (internal_wr_ptr == 11'd883) ) ? wr_data : cam_loc883;
	cam_loc884 <= (internal_wr_en & (internal_wr_ptr == 11'd884) ) ? wr_data : cam_loc884;
	cam_loc885 <= (internal_wr_en & (internal_wr_ptr == 11'd885) ) ? wr_data : cam_loc885;
	cam_loc886 <= (internal_wr_en & (internal_wr_ptr == 11'd886) ) ? wr_data : cam_loc886;
	cam_loc887 <= (internal_wr_en & (internal_wr_ptr == 11'd887) ) ? wr_data : cam_loc887;
	cam_loc888 <= (internal_wr_en & (internal_wr_ptr == 11'd888) ) ? wr_data : cam_loc888;
	cam_loc889 <= (internal_wr_en & (internal_wr_ptr == 11'd889) ) ? wr_data : cam_loc889;
	cam_loc890 <= (internal_wr_en & (internal_wr_ptr == 11'd890) ) ? wr_data : cam_loc890;
	cam_loc891 <= (internal_wr_en & (internal_wr_ptr == 11'd891) ) ? wr_data : cam_loc891;
	cam_loc892 <= (internal_wr_en & (internal_wr_ptr == 11'd892) ) ? wr_data : cam_loc892;
	cam_loc893 <= (internal_wr_en & (internal_wr_ptr == 11'd893) ) ? wr_data : cam_loc893;
	cam_loc894 <= (internal_wr_en & (internal_wr_ptr == 11'd894) ) ? wr_data : cam_loc894;
	cam_loc895 <= (internal_wr_en & (internal_wr_ptr == 11'd895) ) ? wr_data : cam_loc895;
	cam_loc896 <= (internal_wr_en & (internal_wr_ptr == 11'd896) ) ? wr_data : cam_loc896;
	cam_loc897 <= (internal_wr_en & (internal_wr_ptr == 11'd897) ) ? wr_data : cam_loc897;
	cam_loc898 <= (internal_wr_en & (internal_wr_ptr == 11'd898) ) ? wr_data : cam_loc898;
	cam_loc899 <= (internal_wr_en & (internal_wr_ptr == 11'd899) ) ? wr_data : cam_loc899;
	cam_loc900 <= (internal_wr_en & (internal_wr_ptr == 11'd900) ) ? wr_data : cam_loc900;
	cam_loc901 <= (internal_wr_en & (internal_wr_ptr == 11'd901) ) ? wr_data : cam_loc901;
	cam_loc902 <= (internal_wr_en & (internal_wr_ptr == 11'd902) ) ? wr_data : cam_loc902;
	cam_loc903 <= (internal_wr_en & (internal_wr_ptr == 11'd903) ) ? wr_data : cam_loc903;
	cam_loc904 <= (internal_wr_en & (internal_wr_ptr == 11'd904) ) ? wr_data : cam_loc904;
	cam_loc905 <= (internal_wr_en & (internal_wr_ptr == 11'd905) ) ? wr_data : cam_loc905;
	cam_loc906 <= (internal_wr_en & (internal_wr_ptr == 11'd906) ) ? wr_data : cam_loc906;
	cam_loc907 <= (internal_wr_en & (internal_wr_ptr == 11'd907) ) ? wr_data : cam_loc907;
	cam_loc908 <= (internal_wr_en & (internal_wr_ptr == 11'd908) ) ? wr_data : cam_loc908;
	cam_loc909 <= (internal_wr_en & (internal_wr_ptr == 11'd909) ) ? wr_data : cam_loc909;
	cam_loc910 <= (internal_wr_en & (internal_wr_ptr == 11'd910) ) ? wr_data : cam_loc910;
	cam_loc911 <= (internal_wr_en & (internal_wr_ptr == 11'd911) ) ? wr_data : cam_loc911;
	cam_loc912 <= (internal_wr_en & (internal_wr_ptr == 11'd912) ) ? wr_data : cam_loc912;
	cam_loc913 <= (internal_wr_en & (internal_wr_ptr == 11'd913) ) ? wr_data : cam_loc913;
	cam_loc914 <= (internal_wr_en & (internal_wr_ptr == 11'd914) ) ? wr_data : cam_loc914;
	cam_loc915 <= (internal_wr_en & (internal_wr_ptr == 11'd915) ) ? wr_data : cam_loc915;
	cam_loc916 <= (internal_wr_en & (internal_wr_ptr == 11'd916) ) ? wr_data : cam_loc916;
	cam_loc917 <= (internal_wr_en & (internal_wr_ptr == 11'd917) ) ? wr_data : cam_loc917;
	cam_loc918 <= (internal_wr_en & (internal_wr_ptr == 11'd918) ) ? wr_data : cam_loc918;
	cam_loc919 <= (internal_wr_en & (internal_wr_ptr == 11'd919) ) ? wr_data : cam_loc919;
	cam_loc920 <= (internal_wr_en & (internal_wr_ptr == 11'd920) ) ? wr_data : cam_loc920;
	cam_loc921 <= (internal_wr_en & (internal_wr_ptr == 11'd921) ) ? wr_data : cam_loc921;
	cam_loc922 <= (internal_wr_en & (internal_wr_ptr == 11'd922) ) ? wr_data : cam_loc922;
	cam_loc923 <= (internal_wr_en & (internal_wr_ptr == 11'd923) ) ? wr_data : cam_loc923;
	cam_loc924 <= (internal_wr_en & (internal_wr_ptr == 11'd924) ) ? wr_data : cam_loc924;
	cam_loc925 <= (internal_wr_en & (internal_wr_ptr == 11'd925) ) ? wr_data : cam_loc925;
	cam_loc926 <= (internal_wr_en & (internal_wr_ptr == 11'd926) ) ? wr_data : cam_loc926;
	cam_loc927 <= (internal_wr_en & (internal_wr_ptr == 11'd927) ) ? wr_data : cam_loc927;
	cam_loc928 <= (internal_wr_en & (internal_wr_ptr == 11'd928) ) ? wr_data : cam_loc928;
	cam_loc929 <= (internal_wr_en & (internal_wr_ptr == 11'd929) ) ? wr_data : cam_loc929;
	cam_loc930 <= (internal_wr_en & (internal_wr_ptr == 11'd930) ) ? wr_data : cam_loc930;
	cam_loc931 <= (internal_wr_en & (internal_wr_ptr == 11'd931) ) ? wr_data : cam_loc931;
	cam_loc932 <= (internal_wr_en & (internal_wr_ptr == 11'd932) ) ? wr_data : cam_loc932;
	cam_loc933 <= (internal_wr_en & (internal_wr_ptr == 11'd933) ) ? wr_data : cam_loc933;
	cam_loc934 <= (internal_wr_en & (internal_wr_ptr == 11'd934) ) ? wr_data : cam_loc934;
	cam_loc935 <= (internal_wr_en & (internal_wr_ptr == 11'd935) ) ? wr_data : cam_loc935;
	cam_loc936 <= (internal_wr_en & (internal_wr_ptr == 11'd936) ) ? wr_data : cam_loc936;
	cam_loc937 <= (internal_wr_en & (internal_wr_ptr == 11'd937) ) ? wr_data : cam_loc937;
	cam_loc938 <= (internal_wr_en & (internal_wr_ptr == 11'd938) ) ? wr_data : cam_loc938;
	cam_loc939 <= (internal_wr_en & (internal_wr_ptr == 11'd939) ) ? wr_data : cam_loc939;
	cam_loc940 <= (internal_wr_en & (internal_wr_ptr == 11'd940) ) ? wr_data : cam_loc940;
	cam_loc941 <= (internal_wr_en & (internal_wr_ptr == 11'd941) ) ? wr_data : cam_loc941;
	cam_loc942 <= (internal_wr_en & (internal_wr_ptr == 11'd942) ) ? wr_data : cam_loc942;
	cam_loc943 <= (internal_wr_en & (internal_wr_ptr == 11'd943) ) ? wr_data : cam_loc943;
	cam_loc944 <= (internal_wr_en & (internal_wr_ptr == 11'd944) ) ? wr_data : cam_loc944;
	cam_loc945 <= (internal_wr_en & (internal_wr_ptr == 11'd945) ) ? wr_data : cam_loc945;
	cam_loc946 <= (internal_wr_en & (internal_wr_ptr == 11'd946) ) ? wr_data : cam_loc946;
	cam_loc947 <= (internal_wr_en & (internal_wr_ptr == 11'd947) ) ? wr_data : cam_loc947;
	cam_loc948 <= (internal_wr_en & (internal_wr_ptr == 11'd948) ) ? wr_data : cam_loc948;
	cam_loc949 <= (internal_wr_en & (internal_wr_ptr == 11'd949) ) ? wr_data : cam_loc949;
	cam_loc950 <= (internal_wr_en & (internal_wr_ptr == 11'd950) ) ? wr_data : cam_loc950;
	cam_loc951 <= (internal_wr_en & (internal_wr_ptr == 11'd951) ) ? wr_data : cam_loc951;
	cam_loc952 <= (internal_wr_en & (internal_wr_ptr == 11'd952) ) ? wr_data : cam_loc952;
	cam_loc953 <= (internal_wr_en & (internal_wr_ptr == 11'd953) ) ? wr_data : cam_loc953;
	cam_loc954 <= (internal_wr_en & (internal_wr_ptr == 11'd954) ) ? wr_data : cam_loc954;
	cam_loc955 <= (internal_wr_en & (internal_wr_ptr == 11'd955) ) ? wr_data : cam_loc955;
	cam_loc956 <= (internal_wr_en & (internal_wr_ptr == 11'd956) ) ? wr_data : cam_loc956;
	cam_loc957 <= (internal_wr_en & (internal_wr_ptr == 11'd957) ) ? wr_data : cam_loc957;
	cam_loc958 <= (internal_wr_en & (internal_wr_ptr == 11'd958) ) ? wr_data : cam_loc958;
	cam_loc959 <= (internal_wr_en & (internal_wr_ptr == 11'd959) ) ? wr_data : cam_loc959;
	cam_loc960 <= (internal_wr_en & (internal_wr_ptr == 11'd960) ) ? wr_data : cam_loc960;
	cam_loc961 <= (internal_wr_en & (internal_wr_ptr == 11'd961) ) ? wr_data : cam_loc961;
	cam_loc962 <= (internal_wr_en & (internal_wr_ptr == 11'd962) ) ? wr_data : cam_loc962;
	cam_loc963 <= (internal_wr_en & (internal_wr_ptr == 11'd963) ) ? wr_data : cam_loc963;
	cam_loc964 <= (internal_wr_en & (internal_wr_ptr == 11'd964) ) ? wr_data : cam_loc964;
	cam_loc965 <= (internal_wr_en & (internal_wr_ptr == 11'd965) ) ? wr_data : cam_loc965;
	cam_loc966 <= (internal_wr_en & (internal_wr_ptr == 11'd966) ) ? wr_data : cam_loc966;
	cam_loc967 <= (internal_wr_en & (internal_wr_ptr == 11'd967) ) ? wr_data : cam_loc967;
	cam_loc968 <= (internal_wr_en & (internal_wr_ptr == 11'd968) ) ? wr_data : cam_loc968;
	cam_loc969 <= (internal_wr_en & (internal_wr_ptr == 11'd969) ) ? wr_data : cam_loc969;
	cam_loc970 <= (internal_wr_en & (internal_wr_ptr == 11'd970) ) ? wr_data : cam_loc970;
	cam_loc971 <= (internal_wr_en & (internal_wr_ptr == 11'd971) ) ? wr_data : cam_loc971;
	cam_loc972 <= (internal_wr_en & (internal_wr_ptr == 11'd972) ) ? wr_data : cam_loc972;
	cam_loc973 <= (internal_wr_en & (internal_wr_ptr == 11'd973) ) ? wr_data : cam_loc973;
	cam_loc974 <= (internal_wr_en & (internal_wr_ptr == 11'd974) ) ? wr_data : cam_loc974;
	cam_loc975 <= (internal_wr_en & (internal_wr_ptr == 11'd975) ) ? wr_data : cam_loc975;
	cam_loc976 <= (internal_wr_en & (internal_wr_ptr == 11'd976) ) ? wr_data : cam_loc976;
	cam_loc977 <= (internal_wr_en & (internal_wr_ptr == 11'd977) ) ? wr_data : cam_loc977;
	cam_loc978 <= (internal_wr_en & (internal_wr_ptr == 11'd978) ) ? wr_data : cam_loc978;
	cam_loc979 <= (internal_wr_en & (internal_wr_ptr == 11'd979) ) ? wr_data : cam_loc979;
	cam_loc980 <= (internal_wr_en & (internal_wr_ptr == 11'd980) ) ? wr_data : cam_loc980;
	cam_loc981 <= (internal_wr_en & (internal_wr_ptr == 11'd981) ) ? wr_data : cam_loc981;
	cam_loc982 <= (internal_wr_en & (internal_wr_ptr == 11'd982) ) ? wr_data : cam_loc982;
	cam_loc983 <= (internal_wr_en & (internal_wr_ptr == 11'd983) ) ? wr_data : cam_loc983;
	cam_loc984 <= (internal_wr_en & (internal_wr_ptr == 11'd984) ) ? wr_data : cam_loc984;
	cam_loc985 <= (internal_wr_en & (internal_wr_ptr == 11'd985) ) ? wr_data : cam_loc985;
	cam_loc986 <= (internal_wr_en & (internal_wr_ptr == 11'd986) ) ? wr_data : cam_loc986;
	cam_loc987 <= (internal_wr_en & (internal_wr_ptr == 11'd987) ) ? wr_data : cam_loc987;
	cam_loc988 <= (internal_wr_en & (internal_wr_ptr == 11'd988) ) ? wr_data : cam_loc988;
	cam_loc989 <= (internal_wr_en & (internal_wr_ptr == 11'd989) ) ? wr_data : cam_loc989;
	cam_loc990 <= (internal_wr_en & (internal_wr_ptr == 11'd990) ) ? wr_data : cam_loc990;
	cam_loc991 <= (internal_wr_en & (internal_wr_ptr == 11'd991) ) ? wr_data : cam_loc991;
	cam_loc992 <= (internal_wr_en & (internal_wr_ptr == 11'd992) ) ? wr_data : cam_loc992;
	cam_loc993 <= (internal_wr_en & (internal_wr_ptr == 11'd993) ) ? wr_data : cam_loc993;
	cam_loc994 <= (internal_wr_en & (internal_wr_ptr == 11'd994) ) ? wr_data : cam_loc994;
	cam_loc995 <= (internal_wr_en & (internal_wr_ptr == 11'd995) ) ? wr_data : cam_loc995;
	cam_loc996 <= (internal_wr_en & (internal_wr_ptr == 11'd996) ) ? wr_data : cam_loc996;
	cam_loc997 <= (internal_wr_en & (internal_wr_ptr == 11'd997) ) ? wr_data : cam_loc997;
	cam_loc998 <= (internal_wr_en & (internal_wr_ptr == 11'd998) ) ? wr_data : cam_loc998;
	cam_loc999 <= (internal_wr_en & (internal_wr_ptr == 11'd999) ) ? wr_data : cam_loc999;
	cam_loc1000 <= (internal_wr_en & (internal_wr_ptr == 11'd1000) ) ? wr_data : cam_loc1000;
	cam_loc1001 <= (internal_wr_en & (internal_wr_ptr == 11'd1001) ) ? wr_data : cam_loc1001;
	cam_loc1002 <= (internal_wr_en & (internal_wr_ptr == 11'd1002) ) ? wr_data : cam_loc1002;
	cam_loc1003 <= (internal_wr_en & (internal_wr_ptr == 11'd1003) ) ? wr_data : cam_loc1003;
	cam_loc1004 <= (internal_wr_en & (internal_wr_ptr == 11'd1004) ) ? wr_data : cam_loc1004;
	cam_loc1005 <= (internal_wr_en & (internal_wr_ptr == 11'd1005) ) ? wr_data : cam_loc1005;
	cam_loc1006 <= (internal_wr_en & (internal_wr_ptr == 11'd1006) ) ? wr_data : cam_loc1006;
	cam_loc1007 <= (internal_wr_en & (internal_wr_ptr == 11'd1007) ) ? wr_data : cam_loc1007;
	cam_loc1008 <= (internal_wr_en & (internal_wr_ptr == 11'd1008) ) ? wr_data : cam_loc1008;
	cam_loc1009 <= (internal_wr_en & (internal_wr_ptr == 11'd1009) ) ? wr_data : cam_loc1009;
	cam_loc1010 <= (internal_wr_en & (internal_wr_ptr == 11'd1010) ) ? wr_data : cam_loc1010;
	cam_loc1011 <= (internal_wr_en & (internal_wr_ptr == 11'd1011) ) ? wr_data : cam_loc1011;
	cam_loc1012 <= (internal_wr_en & (internal_wr_ptr == 11'd1012) ) ? wr_data : cam_loc1012;
	cam_loc1013 <= (internal_wr_en & (internal_wr_ptr == 11'd1013) ) ? wr_data : cam_loc1013;
	cam_loc1014 <= (internal_wr_en & (internal_wr_ptr == 11'd1014) ) ? wr_data : cam_loc1014;
	cam_loc1015 <= (internal_wr_en & (internal_wr_ptr == 11'd1015) ) ? wr_data : cam_loc1015;
	cam_loc1016 <= (internal_wr_en & (internal_wr_ptr == 11'd1016) ) ? wr_data : cam_loc1016;
	cam_loc1017 <= (internal_wr_en & (internal_wr_ptr == 11'd1017) ) ? wr_data : cam_loc1017;
	cam_loc1018 <= (internal_wr_en & (internal_wr_ptr == 11'd1018) ) ? wr_data : cam_loc1018;
	cam_loc1019 <= (internal_wr_en & (internal_wr_ptr == 11'd1019) ) ? wr_data : cam_loc1019;
	cam_loc1020 <= (internal_wr_en & (internal_wr_ptr == 11'd1020) ) ? wr_data : cam_loc1020;
	cam_loc1021 <= (internal_wr_en & (internal_wr_ptr == 11'd1021) ) ? wr_data : cam_loc1021;
	cam_loc1022 <= (internal_wr_en & (internal_wr_ptr == 11'd1022) ) ? wr_data : cam_loc1022;
	cam_loc1023 <= (internal_wr_en & (internal_wr_ptr == 11'd1023) ) ? wr_data : cam_loc1023;
	cam_loc1024 <= (internal_wr_en & (internal_wr_ptr == 11'd1024) ) ? wr_data : cam_loc1024;
	cam_loc1025 <= (internal_wr_en & (internal_wr_ptr == 11'd1025) ) ? wr_data : cam_loc1025;
	cam_loc1026 <= (internal_wr_en & (internal_wr_ptr == 11'd1026) ) ? wr_data : cam_loc1026;
	cam_loc1027 <= (internal_wr_en & (internal_wr_ptr == 11'd1027) ) ? wr_data : cam_loc1027;
	cam_loc1028 <= (internal_wr_en & (internal_wr_ptr == 11'd1028) ) ? wr_data : cam_loc1028;
	cam_loc1029 <= (internal_wr_en & (internal_wr_ptr == 11'd1029) ) ? wr_data : cam_loc1029;
	cam_loc1030 <= (internal_wr_en & (internal_wr_ptr == 11'd1030) ) ? wr_data : cam_loc1030;
	cam_loc1031 <= (internal_wr_en & (internal_wr_ptr == 11'd1031) ) ? wr_data : cam_loc1031;
	cam_loc1032 <= (internal_wr_en & (internal_wr_ptr == 11'd1032) ) ? wr_data : cam_loc1032;
	cam_loc1033 <= (internal_wr_en & (internal_wr_ptr == 11'd1033) ) ? wr_data : cam_loc1033;
	cam_loc1034 <= (internal_wr_en & (internal_wr_ptr == 11'd1034) ) ? wr_data : cam_loc1034;
	cam_loc1035 <= (internal_wr_en & (internal_wr_ptr == 11'd1035) ) ? wr_data : cam_loc1035;
	cam_loc1036 <= (internal_wr_en & (internal_wr_ptr == 11'd1036) ) ? wr_data : cam_loc1036;
	cam_loc1037 <= (internal_wr_en & (internal_wr_ptr == 11'd1037) ) ? wr_data : cam_loc1037;
	cam_loc1038 <= (internal_wr_en & (internal_wr_ptr == 11'd1038) ) ? wr_data : cam_loc1038;
	cam_loc1039 <= (internal_wr_en & (internal_wr_ptr == 11'd1039) ) ? wr_data : cam_loc1039;
	cam_loc1040 <= (internal_wr_en & (internal_wr_ptr == 11'd1040) ) ? wr_data : cam_loc1040;
	cam_loc1041 <= (internal_wr_en & (internal_wr_ptr == 11'd1041) ) ? wr_data : cam_loc1041;
	cam_loc1042 <= (internal_wr_en & (internal_wr_ptr == 11'd1042) ) ? wr_data : cam_loc1042;
	cam_loc1043 <= (internal_wr_en & (internal_wr_ptr == 11'd1043) ) ? wr_data : cam_loc1043;
	cam_loc1044 <= (internal_wr_en & (internal_wr_ptr == 11'd1044) ) ? wr_data : cam_loc1044;
	cam_loc1045 <= (internal_wr_en & (internal_wr_ptr == 11'd1045) ) ? wr_data : cam_loc1045;
	cam_loc1046 <= (internal_wr_en & (internal_wr_ptr == 11'd1046) ) ? wr_data : cam_loc1046;
	cam_loc1047 <= (internal_wr_en & (internal_wr_ptr == 11'd1047) ) ? wr_data : cam_loc1047;
	cam_loc1048 <= (internal_wr_en & (internal_wr_ptr == 11'd1048) ) ? wr_data : cam_loc1048;
	cam_loc1049 <= (internal_wr_en & (internal_wr_ptr == 11'd1049) ) ? wr_data : cam_loc1049;
	cam_loc1050 <= (internal_wr_en & (internal_wr_ptr == 11'd1050) ) ? wr_data : cam_loc1050;
	cam_loc1051 <= (internal_wr_en & (internal_wr_ptr == 11'd1051) ) ? wr_data : cam_loc1051;
	cam_loc1052 <= (internal_wr_en & (internal_wr_ptr == 11'd1052) ) ? wr_data : cam_loc1052;
	cam_loc1053 <= (internal_wr_en & (internal_wr_ptr == 11'd1053) ) ? wr_data : cam_loc1053;
	cam_loc1054 <= (internal_wr_en & (internal_wr_ptr == 11'd1054) ) ? wr_data : cam_loc1054;
	cam_loc1055 <= (internal_wr_en & (internal_wr_ptr == 11'd1055) ) ? wr_data : cam_loc1055;
	cam_loc1056 <= (internal_wr_en & (internal_wr_ptr == 11'd1056) ) ? wr_data : cam_loc1056;
	cam_loc1057 <= (internal_wr_en & (internal_wr_ptr == 11'd1057) ) ? wr_data : cam_loc1057;
	cam_loc1058 <= (internal_wr_en & (internal_wr_ptr == 11'd1058) ) ? wr_data : cam_loc1058;
	cam_loc1059 <= (internal_wr_en & (internal_wr_ptr == 11'd1059) ) ? wr_data : cam_loc1059;
	cam_loc1060 <= (internal_wr_en & (internal_wr_ptr == 11'd1060) ) ? wr_data : cam_loc1060;
	cam_loc1061 <= (internal_wr_en & (internal_wr_ptr == 11'd1061) ) ? wr_data : cam_loc1061;
	cam_loc1062 <= (internal_wr_en & (internal_wr_ptr == 11'd1062) ) ? wr_data : cam_loc1062;
	cam_loc1063 <= (internal_wr_en & (internal_wr_ptr == 11'd1063) ) ? wr_data : cam_loc1063;
	cam_loc1064 <= (internal_wr_en & (internal_wr_ptr == 11'd1064) ) ? wr_data : cam_loc1064;
	cam_loc1065 <= (internal_wr_en & (internal_wr_ptr == 11'd1065) ) ? wr_data : cam_loc1065;
	cam_loc1066 <= (internal_wr_en & (internal_wr_ptr == 11'd1066) ) ? wr_data : cam_loc1066;
	cam_loc1067 <= (internal_wr_en & (internal_wr_ptr == 11'd1067) ) ? wr_data : cam_loc1067;
	cam_loc1068 <= (internal_wr_en & (internal_wr_ptr == 11'd1068) ) ? wr_data : cam_loc1068;
	cam_loc1069 <= (internal_wr_en & (internal_wr_ptr == 11'd1069) ) ? wr_data : cam_loc1069;
	cam_loc1070 <= (internal_wr_en & (internal_wr_ptr == 11'd1070) ) ? wr_data : cam_loc1070;
	cam_loc1071 <= (internal_wr_en & (internal_wr_ptr == 11'd1071) ) ? wr_data : cam_loc1071;
	cam_loc1072 <= (internal_wr_en & (internal_wr_ptr == 11'd1072) ) ? wr_data : cam_loc1072;
	cam_loc1073 <= (internal_wr_en & (internal_wr_ptr == 11'd1073) ) ? wr_data : cam_loc1073;
	cam_loc1074 <= (internal_wr_en & (internal_wr_ptr == 11'd1074) ) ? wr_data : cam_loc1074;
	cam_loc1075 <= (internal_wr_en & (internal_wr_ptr == 11'd1075) ) ? wr_data : cam_loc1075;
	cam_loc1076 <= (internal_wr_en & (internal_wr_ptr == 11'd1076) ) ? wr_data : cam_loc1076;
	cam_loc1077 <= (internal_wr_en & (internal_wr_ptr == 11'd1077) ) ? wr_data : cam_loc1077;
	cam_loc1078 <= (internal_wr_en & (internal_wr_ptr == 11'd1078) ) ? wr_data : cam_loc1078;
	cam_loc1079 <= (internal_wr_en & (internal_wr_ptr == 11'd1079) ) ? wr_data : cam_loc1079;
	cam_loc1080 <= (internal_wr_en & (internal_wr_ptr == 11'd1080) ) ? wr_data : cam_loc1080;
	cam_loc1081 <= (internal_wr_en & (internal_wr_ptr == 11'd1081) ) ? wr_data : cam_loc1081;
	cam_loc1082 <= (internal_wr_en & (internal_wr_ptr == 11'd1082) ) ? wr_data : cam_loc1082;
	cam_loc1083 <= (internal_wr_en & (internal_wr_ptr == 11'd1083) ) ? wr_data : cam_loc1083;
	cam_loc1084 <= (internal_wr_en & (internal_wr_ptr == 11'd1084) ) ? wr_data : cam_loc1084;
	cam_loc1085 <= (internal_wr_en & (internal_wr_ptr == 11'd1085) ) ? wr_data : cam_loc1085;
	cam_loc1086 <= (internal_wr_en & (internal_wr_ptr == 11'd1086) ) ? wr_data : cam_loc1086;
	cam_loc1087 <= (internal_wr_en & (internal_wr_ptr == 11'd1087) ) ? wr_data : cam_loc1087;
	cam_loc1088 <= (internal_wr_en & (internal_wr_ptr == 11'd1088) ) ? wr_data : cam_loc1088;
	cam_loc1089 <= (internal_wr_en & (internal_wr_ptr == 11'd1089) ) ? wr_data : cam_loc1089;
	cam_loc1090 <= (internal_wr_en & (internal_wr_ptr == 11'd1090) ) ? wr_data : cam_loc1090;
	cam_loc1091 <= (internal_wr_en & (internal_wr_ptr == 11'd1091) ) ? wr_data : cam_loc1091;
	cam_loc1092 <= (internal_wr_en & (internal_wr_ptr == 11'd1092) ) ? wr_data : cam_loc1092;
	cam_loc1093 <= (internal_wr_en & (internal_wr_ptr == 11'd1093) ) ? wr_data : cam_loc1093;
	cam_loc1094 <= (internal_wr_en & (internal_wr_ptr == 11'd1094) ) ? wr_data : cam_loc1094;
	cam_loc1095 <= (internal_wr_en & (internal_wr_ptr == 11'd1095) ) ? wr_data : cam_loc1095;
	cam_loc1096 <= (internal_wr_en & (internal_wr_ptr == 11'd1096) ) ? wr_data : cam_loc1096;
	cam_loc1097 <= (internal_wr_en & (internal_wr_ptr == 11'd1097) ) ? wr_data : cam_loc1097;
	cam_loc1098 <= (internal_wr_en & (internal_wr_ptr == 11'd1098) ) ? wr_data : cam_loc1098;
	cam_loc1099 <= (internal_wr_en & (internal_wr_ptr == 11'd1099) ) ? wr_data : cam_loc1099;


end

wire assign snoop_match = freedup_loc_ready) & (

(snoop_in == cam_loc0[14:0]) |
 (snoop_in == cam_loc1[14:0]) |
 (snoop_in == cam_loc2[14:0]) |
 (snoop_in == cam_loc3[14:0]) |
 (snoop_in == cam_loc4[14:0]) |
 (snoop_in == cam_loc5[14:0]) |
 (snoop_in == cam_loc6[14:0]) |
 (snoop_in == cam_loc7[14:0]) |
 (snoop_in == cam_loc8[14:0]) |
 (snoop_in == cam_loc9[14:0]) |
 (snoop_in == cam_loc10[14:0]) |
 (snoop_in == cam_loc11[14:0]) |
 (snoop_in == cam_loc12[14:0]) |
 (snoop_in == cam_loc13[14:0]) |
 (snoop_in == cam_loc14[14:0]) |
 (snoop_in == cam_loc15[14:0]) |
 (snoop_in == cam_loc16[14:0]) |
 (snoop_in == cam_loc17[14:0]) |
 (snoop_in == cam_loc18[14:0]) |
 (snoop_in == cam_loc19[14:0]) |
 (snoop_in == cam_loc20[14:0]) |
 (snoop_in == cam_loc21[14:0]) |
 (snoop_in == cam_loc22[14:0]) |
 (snoop_in == cam_loc23[14:0]) |
 (snoop_in == cam_loc24[14:0]) |
 (snoop_in == cam_loc25[14:0]) |
 (snoop_in == cam_loc26[14:0]) |
 (snoop_in == cam_loc27[14:0]) |
 (snoop_in == cam_loc28[14:0]) |
 (snoop_in == cam_loc29[14:0]) |
 (snoop_in == cam_loc30[14:0]) |
 (snoop_in == cam_loc31[14:0]) |
 (snoop_in == cam_loc32[14:0]) |
 (snoop_in == cam_loc33[14:0]) |
 (snoop_in == cam_loc34[14:0]) |
 (snoop_in == cam_loc35[14:0]) |
 (snoop_in == cam_loc36[14:0]) |
 (snoop_in == cam_loc37[14:0]) |
 (snoop_in == cam_loc38[14:0]) |
 (snoop_in == cam_loc39[14:0]) |
 (snoop_in == cam_loc40[14:0]) |
 (snoop_in == cam_loc41[14:0]) |
 (snoop_in == cam_loc42[14:0]) |
 (snoop_in == cam_loc43[14:0]) |
 (snoop_in == cam_loc44[14:0]) |
 (snoop_in == cam_loc45[14:0]) |
 (snoop_in == cam_loc46[14:0]) |
 (snoop_in == cam_loc47[14:0]) |
 (snoop_in == cam_loc48[14:0]) |
 (snoop_in == cam_loc49[14:0]) |
 (snoop_in == cam_loc50[14:0]) |
 (snoop_in == cam_loc51[14:0]) |
 (snoop_in == cam_loc52[14:0]) |
 (snoop_in == cam_loc53[14:0]) |
 (snoop_in == cam_loc54[14:0]) |
 (snoop_in == cam_loc55[14:0]) |
 (snoop_in == cam_loc56[14:0]) |
 (snoop_in == cam_loc57[14:0]) |
 (snoop_in == cam_loc58[14:0]) |
 (snoop_in == cam_loc59[14:0]) |
 (snoop_in == cam_loc60[14:0]) |
 (snoop_in == cam_loc61[14:0]) |
 (snoop_in == cam_loc62[14:0]) |
 (snoop_in == cam_loc63[14:0]) |
 (snoop_in == cam_loc64[14:0]) |
 (snoop_in == cam_loc65[14:0]) |
 (snoop_in == cam_loc66[14:0]) |
 (snoop_in == cam_loc67[14:0]) |
 (snoop_in == cam_loc68[14:0]) |
 (snoop_in == cam_loc69[14:0]) |
 (snoop_in == cam_loc70[14:0]) |
 (snoop_in == cam_loc71[14:0]) |
 (snoop_in == cam_loc72[14:0]) |
 (snoop_in == cam_loc73[14:0]) |
 (snoop_in == cam_loc74[14:0]) |
 (snoop_in == cam_loc75[14:0]) |
 (snoop_in == cam_loc76[14:0]) |
 (snoop_in == cam_loc77[14:0]) |
 (snoop_in == cam_loc78[14:0]) |
 (snoop_in == cam_loc79[14:0]) |
 (snoop_in == cam_loc80[14:0]) |
 (snoop_in == cam_loc81[14:0]) |
 (snoop_in == cam_loc82[14:0]) |
 (snoop_in == cam_loc83[14:0]) |
 (snoop_in == cam_loc84[14:0]) |
 (snoop_in == cam_loc85[14:0]) |
 (snoop_in == cam_loc86[14:0]) |
 (snoop_in == cam_loc87[14:0]) |
 (snoop_in == cam_loc88[14:0]) |
 (snoop_in == cam_loc89[14:0]) |
 (snoop_in == cam_loc90[14:0]) |
 (snoop_in == cam_loc91[14:0]) |
 (snoop_in == cam_loc92[14:0]) |
 (snoop_in == cam_loc93[14:0]) |
 (snoop_in == cam_loc94[14:0]) |
 (snoop_in == cam_loc95[14:0]) |
 (snoop_in == cam_loc96[14:0]) |
 (snoop_in == cam_loc97[14:0]) |
 (snoop_in == cam_loc98[14:0]) |
 (snoop_in == cam_loc99[14:0]) |
 (snoop_in == cam_loc100[14:0]) |
 (snoop_in == cam_loc101[14:0]) |
 (snoop_in == cam_loc102[14:0]) |
 (snoop_in == cam_loc103[14:0]) |
 (snoop_in == cam_loc104[14:0]) |
 (snoop_in == cam_loc105[14:0]) |
 (snoop_in == cam_loc106[14:0]) |
 (snoop_in == cam_loc107[14:0]) |
 (snoop_in == cam_loc108[14:0]) |
 (snoop_in == cam_loc109[14:0]) |
 (snoop_in == cam_loc110[14:0]) |
 (snoop_in == cam_loc111[14:0]) |
 (snoop_in == cam_loc112[14:0]) |
 (snoop_in == cam_loc113[14:0]) |
 (snoop_in == cam_loc114[14:0]) |
 (snoop_in == cam_loc115[14:0]) |
 (snoop_in == cam_loc116[14:0]) |
 (snoop_in == cam_loc117[14:0]) |
 (snoop_in == cam_loc118[14:0]) |
 (snoop_in == cam_loc119[14:0]) |
 (snoop_in == cam_loc120[14:0]) |
 (snoop_in == cam_loc121[14:0]) |
 (snoop_in == cam_loc122[14:0]) |
 (snoop_in == cam_loc123[14:0]) |
 (snoop_in == cam_loc124[14:0]) |
 (snoop_in == cam_loc125[14:0]) |
 (snoop_in == cam_loc126[14:0]) |
 (snoop_in == cam_loc127[14:0]) |
 (snoop_in == cam_loc128[14:0]) |
 (snoop_in == cam_loc129[14:0]) |
 (snoop_in == cam_loc130[14:0]) |
 (snoop_in == cam_loc131[14:0]) |
 (snoop_in == cam_loc132[14:0]) |
 (snoop_in == cam_loc133[14:0]) |
 (snoop_in == cam_loc134[14:0]) |
 (snoop_in == cam_loc135[14:0]) |
 (snoop_in == cam_loc136[14:0]) |
 (snoop_in == cam_loc137[14:0]) |
 (snoop_in == cam_loc138[14:0]) |
 (snoop_in == cam_loc139[14:0]) |
 (snoop_in == cam_loc140[14:0]) |
 (snoop_in == cam_loc141[14:0]) |
 (snoop_in == cam_loc142[14:0]) |
 (snoop_in == cam_loc143[14:0]) |
 (snoop_in == cam_loc144[14:0]) |
 (snoop_in == cam_loc145[14:0]) |
 (snoop_in == cam_loc146[14:0]) |
 (snoop_in == cam_loc147[14:0]) |
 (snoop_in == cam_loc148[14:0]) |
 (snoop_in == cam_loc149[14:0]) |
 (snoop_in == cam_loc150[14:0]) |
 (snoop_in == cam_loc151[14:0]) |
 (snoop_in == cam_loc152[14:0]) |
 (snoop_in == cam_loc153[14:0]) |
 (snoop_in == cam_loc154[14:0]) |
 (snoop_in == cam_loc155[14:0]) |
 (snoop_in == cam_loc156[14:0]) |
 (snoop_in == cam_loc157[14:0]) |
 (snoop_in == cam_loc158[14:0]) |
 (snoop_in == cam_loc159[14:0]) |
 (snoop_in == cam_loc160[14:0]) |
 (snoop_in == cam_loc161[14:0]) |
 (snoop_in == cam_loc162[14:0]) |
 (snoop_in == cam_loc163[14:0]) |
 (snoop_in == cam_loc164[14:0]) |
 (snoop_in == cam_loc165[14:0]) |
 (snoop_in == cam_loc166[14:0]) |
 (snoop_in == cam_loc167[14:0]) |
 (snoop_in == cam_loc168[14:0]) |
 (snoop_in == cam_loc169[14:0]) |
 (snoop_in == cam_loc170[14:0]) |
 (snoop_in == cam_loc171[14:0]) |
 (snoop_in == cam_loc172[14:0]) |
 (snoop_in == cam_loc173[14:0]) |
 (snoop_in == cam_loc174[14:0]) |
 (snoop_in == cam_loc175[14:0]) |
 (snoop_in == cam_loc176[14:0]) |
 (snoop_in == cam_loc177[14:0]) |
 (snoop_in == cam_loc178[14:0]) |
 (snoop_in == cam_loc179[14:0]) |
 (snoop_in == cam_loc180[14:0]) |
 (snoop_in == cam_loc181[14:0]) |
 (snoop_in == cam_loc182[14:0]) |
 (snoop_in == cam_loc183[14:0]) |
 (snoop_in == cam_loc184[14:0]) |
 (snoop_in == cam_loc185[14:0]) |
 (snoop_in == cam_loc186[14:0]) |
 (snoop_in == cam_loc187[14:0]) |
 (snoop_in == cam_loc188[14:0]) |
 (snoop_in == cam_loc189[14:0]) |
 (snoop_in == cam_loc190[14:0]) |
 (snoop_in == cam_loc191[14:0]) |
 (snoop_in == cam_loc192[14:0]) |
 (snoop_in == cam_loc193[14:0]) |
 (snoop_in == cam_loc194[14:0]) |
 (snoop_in == cam_loc195[14:0]) |
 (snoop_in == cam_loc196[14:0]) |
 (snoop_in == cam_loc197[14:0]) |
 (snoop_in == cam_loc198[14:0]) |
 (snoop_in == cam_loc199[14:0]) |
 (snoop_in == cam_loc200[14:0]) |
 (snoop_in == cam_loc201[14:0]) |
 (snoop_in == cam_loc202[14:0]) |
 (snoop_in == cam_loc203[14:0]) |
 (snoop_in == cam_loc204[14:0]) |
 (snoop_in == cam_loc205[14:0]) |
 (snoop_in == cam_loc206[14:0]) |
 (snoop_in == cam_loc207[14:0]) |
 (snoop_in == cam_loc208[14:0]) |
 (snoop_in == cam_loc209[14:0]) |
 (snoop_in == cam_loc210[14:0]) |
 (snoop_in == cam_loc211[14:0]) |
 (snoop_in == cam_loc212[14:0]) |
 (snoop_in == cam_loc213[14:0]) |
 (snoop_in == cam_loc214[14:0]) |
 (snoop_in == cam_loc215[14:0]) |
 (snoop_in == cam_loc216[14:0]) |
 (snoop_in == cam_loc217[14:0]) |
 (snoop_in == cam_loc218[14:0]) |
 (snoop_in == cam_loc219[14:0]) |
 (snoop_in == cam_loc220[14:0]) |
 (snoop_in == cam_loc221[14:0]) |
 (snoop_in == cam_loc222[14:0]) |
 (snoop_in == cam_loc223[14:0]) |
 (snoop_in == cam_loc224[14:0]) |
 (snoop_in == cam_loc225[14:0]) |
 (snoop_in == cam_loc226[14:0]) |
 (snoop_in == cam_loc227[14:0]) |
 (snoop_in == cam_loc228[14:0]) |
 (snoop_in == cam_loc229[14:0]) |
 (snoop_in == cam_loc230[14:0]) |
 (snoop_in == cam_loc231[14:0]) |
 (snoop_in == cam_loc232[14:0]) |
 (snoop_in == cam_loc233[14:0]) |
 (snoop_in == cam_loc234[14:0]) |
 (snoop_in == cam_loc235[14:0]) |
 (snoop_in == cam_loc236[14:0]) |
 (snoop_in == cam_loc237[14:0]) |
 (snoop_in == cam_loc238[14:0]) |
 (snoop_in == cam_loc239[14:0]) |
 (snoop_in == cam_loc240[14:0]) |
 (snoop_in == cam_loc241[14:0]) |
 (snoop_in == cam_loc242[14:0]) |
 (snoop_in == cam_loc243[14:0]) |
 (snoop_in == cam_loc244[14:0]) |
 (snoop_in == cam_loc245[14:0]) |
 (snoop_in == cam_loc246[14:0]) |
 (snoop_in == cam_loc247[14:0]) |
 (snoop_in == cam_loc248[14:0]) |
 (snoop_in == cam_loc249[14:0]) |
 (snoop_in == cam_loc250[14:0]) |
 (snoop_in == cam_loc251[14:0]) |
 (snoop_in == cam_loc252[14:0]) |
 (snoop_in == cam_loc253[14:0]) |
 (snoop_in == cam_loc254[14:0]) |
 (snoop_in == cam_loc255[14:0]) |
 (snoop_in == cam_loc256[14:0]) |
 (snoop_in == cam_loc257[14:0]) |
 (snoop_in == cam_loc258[14:0]) |
 (snoop_in == cam_loc259[14:0]) |
 (snoop_in == cam_loc260[14:0]) |
 (snoop_in == cam_loc261[14:0]) |
 (snoop_in == cam_loc262[14:0]) |
 (snoop_in == cam_loc263[14:0]) |
 (snoop_in == cam_loc264[14:0]) |
 (snoop_in == cam_loc265[14:0]) |
 (snoop_in == cam_loc266[14:0]) |
 (snoop_in == cam_loc267[14:0]) |
 (snoop_in == cam_loc268[14:0]) |
 (snoop_in == cam_loc269[14:0]) |
 (snoop_in == cam_loc270[14:0]) |
 (snoop_in == cam_loc271[14:0]) |
 (snoop_in == cam_loc272[14:0]) |
 (snoop_in == cam_loc273[14:0]) |
 (snoop_in == cam_loc274[14:0]) |
 (snoop_in == cam_loc275[14:0]) |
 (snoop_in == cam_loc276[14:0]) |
 (snoop_in == cam_loc277[14:0]) |
 (snoop_in == cam_loc278[14:0]) |
 (snoop_in == cam_loc279[14:0]) |
 (snoop_in == cam_loc280[14:0]) |
 (snoop_in == cam_loc281[14:0]) |
 (snoop_in == cam_loc282[14:0]) |
 (snoop_in == cam_loc283[14:0]) |
 (snoop_in == cam_loc284[14:0]) |
 (snoop_in == cam_loc285[14:0]) |
 (snoop_in == cam_loc286[14:0]) |
 (snoop_in == cam_loc287[14:0]) |
 (snoop_in == cam_loc288[14:0]) |
 (snoop_in == cam_loc289[14:0]) |
 (snoop_in == cam_loc290[14:0]) |
 (snoop_in == cam_loc291[14:0]) |
 (snoop_in == cam_loc292[14:0]) |
 (snoop_in == cam_loc293[14:0]) |
 (snoop_in == cam_loc294[14:0]) |
 (snoop_in == cam_loc295[14:0]) |
 (snoop_in == cam_loc296[14:0]) |
 (snoop_in == cam_loc297[14:0]) |
 (snoop_in == cam_loc298[14:0]) |
 (snoop_in == cam_loc299[14:0]) |
 (snoop_in == cam_loc300[14:0]) |
 (snoop_in == cam_loc301[14:0]) |
 (snoop_in == cam_loc302[14:0]) |
 (snoop_in == cam_loc303[14:0]) |
 (snoop_in == cam_loc304[14:0]) |
 (snoop_in == cam_loc305[14:0]) |
 (snoop_in == cam_loc306[14:0]) |
 (snoop_in == cam_loc307[14:0]) |
 (snoop_in == cam_loc308[14:0]) |
 (snoop_in == cam_loc309[14:0]) |
 (snoop_in == cam_loc310[14:0]) |
 (snoop_in == cam_loc311[14:0]) |
 (snoop_in == cam_loc312[14:0]) |
 (snoop_in == cam_loc313[14:0]) |
 (snoop_in == cam_loc314[14:0]) |
 (snoop_in == cam_loc315[14:0]) |
 (snoop_in == cam_loc316[14:0]) |
 (snoop_in == cam_loc317[14:0]) |
 (snoop_in == cam_loc318[14:0]) |
 (snoop_in == cam_loc319[14:0]) |
 (snoop_in == cam_loc320[14:0]) |
 (snoop_in == cam_loc321[14:0]) |
 (snoop_in == cam_loc322[14:0]) |
 (snoop_in == cam_loc323[14:0]) |
 (snoop_in == cam_loc324[14:0]) |
 (snoop_in == cam_loc325[14:0]) |
 (snoop_in == cam_loc326[14:0]) |
 (snoop_in == cam_loc327[14:0]) |
 (snoop_in == cam_loc328[14:0]) |
 (snoop_in == cam_loc329[14:0]) |
 (snoop_in == cam_loc330[14:0]) |
 (snoop_in == cam_loc331[14:0]) |
 (snoop_in == cam_loc332[14:0]) |
 (snoop_in == cam_loc333[14:0]) |
 (snoop_in == cam_loc334[14:0]) |
 (snoop_in == cam_loc335[14:0]) |
 (snoop_in == cam_loc336[14:0]) |
 (snoop_in == cam_loc337[14:0]) |
 (snoop_in == cam_loc338[14:0]) |
 (snoop_in == cam_loc339[14:0]) |
 (snoop_in == cam_loc340[14:0]) |
 (snoop_in == cam_loc341[14:0]) |
 (snoop_in == cam_loc342[14:0]) |
 (snoop_in == cam_loc343[14:0]) |
 (snoop_in == cam_loc344[14:0]) |
 (snoop_in == cam_loc345[14:0]) |
 (snoop_in == cam_loc346[14:0]) |
 (snoop_in == cam_loc347[14:0]) |
 (snoop_in == cam_loc348[14:0]) |
 (snoop_in == cam_loc349[14:0]) |
 (snoop_in == cam_loc350[14:0]) |
 (snoop_in == cam_loc351[14:0]) |
 (snoop_in == cam_loc352[14:0]) |
 (snoop_in == cam_loc353[14:0]) |
 (snoop_in == cam_loc354[14:0]) |
 (snoop_in == cam_loc355[14:0]) |
 (snoop_in == cam_loc356[14:0]) |
 (snoop_in == cam_loc357[14:0]) |
 (snoop_in == cam_loc358[14:0]) |
 (snoop_in == cam_loc359[14:0]) |
 (snoop_in == cam_loc360[14:0]) |
 (snoop_in == cam_loc361[14:0]) |
 (snoop_in == cam_loc362[14:0]) |
 (snoop_in == cam_loc363[14:0]) |
 (snoop_in == cam_loc364[14:0]) |
 (snoop_in == cam_loc365[14:0]) |
 (snoop_in == cam_loc366[14:0]) |
 (snoop_in == cam_loc367[14:0]) |
 (snoop_in == cam_loc368[14:0]) |
 (snoop_in == cam_loc369[14:0]) |
 (snoop_in == cam_loc370[14:0]) |
 (snoop_in == cam_loc371[14:0]) |
 (snoop_in == cam_loc372[14:0]) |
 (snoop_in == cam_loc373[14:0]) |
 (snoop_in == cam_loc374[14:0]) |
 (snoop_in == cam_loc375[14:0]) |
 (snoop_in == cam_loc376[14:0]) |
 (snoop_in == cam_loc377[14:0]) |
 (snoop_in == cam_loc378[14:0]) |
 (snoop_in == cam_loc379[14:0]) |
 (snoop_in == cam_loc380[14:0]) |
 (snoop_in == cam_loc381[14:0]) |
 (snoop_in == cam_loc382[14:0]) |
 (snoop_in == cam_loc383[14:0]) |
 (snoop_in == cam_loc384[14:0]) |
 (snoop_in == cam_loc385[14:0]) |
 (snoop_in == cam_loc386[14:0]) |
 (snoop_in == cam_loc387[14:0]) |
 (snoop_in == cam_loc388[14:0]) |
 (snoop_in == cam_loc389[14:0]) |
 (snoop_in == cam_loc390[14:0]) |
 (snoop_in == cam_loc391[14:0]) |
 (snoop_in == cam_loc392[14:0]) |
 (snoop_in == cam_loc393[14:0]) |
 (snoop_in == cam_loc394[14:0]) |
 (snoop_in == cam_loc395[14:0]) |
 (snoop_in == cam_loc396[14:0]) |
 (snoop_in == cam_loc397[14:0]) |
 (snoop_in == cam_loc398[14:0]) |
 (snoop_in == cam_loc399[14:0]) |
 (snoop_in == cam_loc400[14:0]) |
 (snoop_in == cam_loc401[14:0]) |
 (snoop_in == cam_loc402[14:0]) |
 (snoop_in == cam_loc403[14:0]) |
 (snoop_in == cam_loc404[14:0]) |
 (snoop_in == cam_loc405[14:0]) |
 (snoop_in == cam_loc406[14:0]) |
 (snoop_in == cam_loc407[14:0]) |
 (snoop_in == cam_loc408[14:0]) |
 (snoop_in == cam_loc409[14:0]) |
 (snoop_in == cam_loc410[14:0]) |
 (snoop_in == cam_loc411[14:0]) |
 (snoop_in == cam_loc412[14:0]) |
 (snoop_in == cam_loc413[14:0]) |
 (snoop_in == cam_loc414[14:0]) |
 (snoop_in == cam_loc415[14:0]) |
 (snoop_in == cam_loc416[14:0]) |
 (snoop_in == cam_loc417[14:0]) |
 (snoop_in == cam_loc418[14:0]) |
 (snoop_in == cam_loc419[14:0]) |
 (snoop_in == cam_loc420[14:0]) |
 (snoop_in == cam_loc421[14:0]) |
 (snoop_in == cam_loc422[14:0]) |
 (snoop_in == cam_loc423[14:0]) |
 (snoop_in == cam_loc424[14:0]) |
 (snoop_in == cam_loc425[14:0]) |
 (snoop_in == cam_loc426[14:0]) |
 (snoop_in == cam_loc427[14:0]) |
 (snoop_in == cam_loc428[14:0]) |
 (snoop_in == cam_loc429[14:0]) |
 (snoop_in == cam_loc430[14:0]) |
 (snoop_in == cam_loc431[14:0]) |
 (snoop_in == cam_loc432[14:0]) |
 (snoop_in == cam_loc433[14:0]) |
 (snoop_in == cam_loc434[14:0]) |
 (snoop_in == cam_loc435[14:0]) |
 (snoop_in == cam_loc436[14:0]) |
 (snoop_in == cam_loc437[14:0]) |
 (snoop_in == cam_loc438[14:0]) |
 (snoop_in == cam_loc439[14:0]) |
 (snoop_in == cam_loc440[14:0]) |
 (snoop_in == cam_loc441[14:0]) |
 (snoop_in == cam_loc442[14:0]) |
 (snoop_in == cam_loc443[14:0]) |
 (snoop_in == cam_loc444[14:0]) |
 (snoop_in == cam_loc445[14:0]) |
 (snoop_in == cam_loc446[14:0]) |
 (snoop_in == cam_loc447[14:0]) |
 (snoop_in == cam_loc448[14:0]) |
 (snoop_in == cam_loc449[14:0]) |
 (snoop_in == cam_loc450[14:0]) |
 (snoop_in == cam_loc451[14:0]) |
 (snoop_in == cam_loc452[14:0]) |
 (snoop_in == cam_loc453[14:0]) |
 (snoop_in == cam_loc454[14:0]) |
 (snoop_in == cam_loc455[14:0]) |
 (snoop_in == cam_loc456[14:0]) |
 (snoop_in == cam_loc457[14:0]) |
 (snoop_in == cam_loc458[14:0]) |
 (snoop_in == cam_loc459[14:0]) |
 (snoop_in == cam_loc460[14:0]) |
 (snoop_in == cam_loc461[14:0]) |
 (snoop_in == cam_loc462[14:0]) |
 (snoop_in == cam_loc463[14:0]) |
 (snoop_in == cam_loc464[14:0]) |
 (snoop_in == cam_loc465[14:0]) |
 (snoop_in == cam_loc466[14:0]) |
 (snoop_in == cam_loc467[14:0]) |
 (snoop_in == cam_loc468[14:0]) |
 (snoop_in == cam_loc469[14:0]) |
 (snoop_in == cam_loc470[14:0]) |
 (snoop_in == cam_loc471[14:0]) |
 (snoop_in == cam_loc472[14:0]) |
 (snoop_in == cam_loc473[14:0]) |
 (snoop_in == cam_loc474[14:0]) |
 (snoop_in == cam_loc475[14:0]) |
 (snoop_in == cam_loc476[14:0]) |
 (snoop_in == cam_loc477[14:0]) |
 (snoop_in == cam_loc478[14:0]) |
 (snoop_in == cam_loc479[14:0]) |
 (snoop_in == cam_loc480[14:0]) |
 (snoop_in == cam_loc481[14:0]) |
 (snoop_in == cam_loc482[14:0]) |
 (snoop_in == cam_loc483[14:0]) |
 (snoop_in == cam_loc484[14:0]) |
 (snoop_in == cam_loc485[14:0]) |
 (snoop_in == cam_loc486[14:0]) |
 (snoop_in == cam_loc487[14:0]) |
 (snoop_in == cam_loc488[14:0]) |
 (snoop_in == cam_loc489[14:0]) |
 (snoop_in == cam_loc490[14:0]) |
 (snoop_in == cam_loc491[14:0]) |
 (snoop_in == cam_loc492[14:0]) |
 (snoop_in == cam_loc493[14:0]) |
 (snoop_in == cam_loc494[14:0]) |
 (snoop_in == cam_loc495[14:0]) |
 (snoop_in == cam_loc496[14:0]) |
 (snoop_in == cam_loc497[14:0]) |
 (snoop_in == cam_loc498[14:0]) |
 (snoop_in == cam_loc499[14:0]) |
 (snoop_in == cam_loc500[14:0]) |
 (snoop_in == cam_loc501[14:0]) |
 (snoop_in == cam_loc502[14:0]) |
 (snoop_in == cam_loc503[14:0]) |
 (snoop_in == cam_loc504[14:0]) |
 (snoop_in == cam_loc505[14:0]) |
 (snoop_in == cam_loc506[14:0]) |
 (snoop_in == cam_loc507[14:0]) |
 (snoop_in == cam_loc508[14:0]) |
 (snoop_in == cam_loc509[14:0]) |
 (snoop_in == cam_loc510[14:0]) |
 (snoop_in == cam_loc511[14:0]) |
 (snoop_in == cam_loc512[14:0]) |
 (snoop_in == cam_loc513[14:0]) |
 (snoop_in == cam_loc514[14:0]) |
 (snoop_in == cam_loc515[14:0]) |
 (snoop_in == cam_loc516[14:0]) |
 (snoop_in == cam_loc517[14:0]) |
 (snoop_in == cam_loc518[14:0]) |
 (snoop_in == cam_loc519[14:0]) |
 (snoop_in == cam_loc520[14:0]) |
 (snoop_in == cam_loc521[14:0]) |
 (snoop_in == cam_loc522[14:0]) |
 (snoop_in == cam_loc523[14:0]) |
 (snoop_in == cam_loc524[14:0]) |
 (snoop_in == cam_loc525[14:0]) |
 (snoop_in == cam_loc526[14:0]) |
 (snoop_in == cam_loc527[14:0]) |
 (snoop_in == cam_loc528[14:0]) |
 (snoop_in == cam_loc529[14:0]) |
 (snoop_in == cam_loc530[14:0]) |
 (snoop_in == cam_loc531[14:0]) |
 (snoop_in == cam_loc532[14:0]) |
 (snoop_in == cam_loc533[14:0]) |
 (snoop_in == cam_loc534[14:0]) |
 (snoop_in == cam_loc535[14:0]) |
 (snoop_in == cam_loc536[14:0]) |
 (snoop_in == cam_loc537[14:0]) |
 (snoop_in == cam_loc538[14:0]) |
 (snoop_in == cam_loc539[14:0]) |
 (snoop_in == cam_loc540[14:0]) |
 (snoop_in == cam_loc541[14:0]) |
 (snoop_in == cam_loc542[14:0]) |
 (snoop_in == cam_loc543[14:0]) |
 (snoop_in == cam_loc544[14:0]) |
 (snoop_in == cam_loc545[14:0]) |
 (snoop_in == cam_loc546[14:0]) |
 (snoop_in == cam_loc547[14:0]) |
 (snoop_in == cam_loc548[14:0]) |
 (snoop_in == cam_loc549[14:0]) |
 (snoop_in == cam_loc550[14:0]) |
 (snoop_in == cam_loc551[14:0]) |
 (snoop_in == cam_loc552[14:0]) |
 (snoop_in == cam_loc553[14:0]) |
 (snoop_in == cam_loc554[14:0]) |
 (snoop_in == cam_loc555[14:0]) |
 (snoop_in == cam_loc556[14:0]) |
 (snoop_in == cam_loc557[14:0]) |
 (snoop_in == cam_loc558[14:0]) |
 (snoop_in == cam_loc559[14:0]) |
 (snoop_in == cam_loc560[14:0]) |
 (snoop_in == cam_loc561[14:0]) |
 (snoop_in == cam_loc562[14:0]) |
 (snoop_in == cam_loc563[14:0]) |
 (snoop_in == cam_loc564[14:0]) |
 (snoop_in == cam_loc565[14:0]) |
 (snoop_in == cam_loc566[14:0]) |
 (snoop_in == cam_loc567[14:0]) |
 (snoop_in == cam_loc568[14:0]) |
 (snoop_in == cam_loc569[14:0]) |
 (snoop_in == cam_loc570[14:0]) |
 (snoop_in == cam_loc571[14:0]) |
 (snoop_in == cam_loc572[14:0]) |
 (snoop_in == cam_loc573[14:0]) |
 (snoop_in == cam_loc574[14:0]) |
 (snoop_in == cam_loc575[14:0]) |
 (snoop_in == cam_loc576[14:0]) |
 (snoop_in == cam_loc577[14:0]) |
 (snoop_in == cam_loc578[14:0]) |
 (snoop_in == cam_loc579[14:0]) |
 (snoop_in == cam_loc580[14:0]) |
 (snoop_in == cam_loc581[14:0]) |
 (snoop_in == cam_loc582[14:0]) |
 (snoop_in == cam_loc583[14:0]) |
 (snoop_in == cam_loc584[14:0]) |
 (snoop_in == cam_loc585[14:0]) |
 (snoop_in == cam_loc586[14:0]) |
 (snoop_in == cam_loc587[14:0]) |
 (snoop_in == cam_loc588[14:0]) |
 (snoop_in == cam_loc589[14:0]) |
 (snoop_in == cam_loc590[14:0]) |
 (snoop_in == cam_loc591[14:0]) |
 (snoop_in == cam_loc592[14:0]) |
 (snoop_in == cam_loc593[14:0]) |
 (snoop_in == cam_loc594[14:0]) |
 (snoop_in == cam_loc595[14:0]) |
 (snoop_in == cam_loc596[14:0]) |
 (snoop_in == cam_loc597[14:0]) |
 (snoop_in == cam_loc598[14:0]) |
 (snoop_in == cam_loc599[14:0]) |
 (snoop_in == cam_loc600[14:0]) |
 (snoop_in == cam_loc601[14:0]) |
 (snoop_in == cam_loc602[14:0]) |
 (snoop_in == cam_loc603[14:0]) |
 (snoop_in == cam_loc604[14:0]) |
 (snoop_in == cam_loc605[14:0]) |
 (snoop_in == cam_loc606[14:0]) |
 (snoop_in == cam_loc607[14:0]) |
 (snoop_in == cam_loc608[14:0]) |
 (snoop_in == cam_loc609[14:0]) |
 (snoop_in == cam_loc610[14:0]) |
 (snoop_in == cam_loc611[14:0]) |
 (snoop_in == cam_loc612[14:0]) |
 (snoop_in == cam_loc613[14:0]) |
 (snoop_in == cam_loc614[14:0]) |
 (snoop_in == cam_loc615[14:0]) |
 (snoop_in == cam_loc616[14:0]) |
 (snoop_in == cam_loc617[14:0]) |
 (snoop_in == cam_loc618[14:0]) |
 (snoop_in == cam_loc619[14:0]) |
 (snoop_in == cam_loc620[14:0]) |
 (snoop_in == cam_loc621[14:0]) |
 (snoop_in == cam_loc622[14:0]) |
 (snoop_in == cam_loc623[14:0]) |
 (snoop_in == cam_loc624[14:0]) |
 (snoop_in == cam_loc625[14:0]) |
 (snoop_in == cam_loc626[14:0]) |
 (snoop_in == cam_loc627[14:0]) |
 (snoop_in == cam_loc628[14:0]) |
 (snoop_in == cam_loc629[14:0]) |
 (snoop_in == cam_loc630[14:0]) |
 (snoop_in == cam_loc631[14:0]) |
 (snoop_in == cam_loc632[14:0]) |
 (snoop_in == cam_loc633[14:0]) |
 (snoop_in == cam_loc634[14:0]) |
 (snoop_in == cam_loc635[14:0]) |
 (snoop_in == cam_loc636[14:0]) |
 (snoop_in == cam_loc637[14:0]) |
 (snoop_in == cam_loc638[14:0]) |
 (snoop_in == cam_loc639[14:0]) |
 (snoop_in == cam_loc640[14:0]) |
 (snoop_in == cam_loc641[14:0]) |
 (snoop_in == cam_loc642[14:0]) |
 (snoop_in == cam_loc643[14:0]) |
 (snoop_in == cam_loc644[14:0]) |
 (snoop_in == cam_loc645[14:0]) |
 (snoop_in == cam_loc646[14:0]) |
 (snoop_in == cam_loc647[14:0]) |
 (snoop_in == cam_loc648[14:0]) |
 (snoop_in == cam_loc649[14:0]) |
 (snoop_in == cam_loc650[14:0]) |
 (snoop_in == cam_loc651[14:0]) |
 (snoop_in == cam_loc652[14:0]) |
 (snoop_in == cam_loc653[14:0]) |
 (snoop_in == cam_loc654[14:0]) |
 (snoop_in == cam_loc655[14:0]) |
 (snoop_in == cam_loc656[14:0]) |
 (snoop_in == cam_loc657[14:0]) |
 (snoop_in == cam_loc658[14:0]) |
 (snoop_in == cam_loc659[14:0]) |
 (snoop_in == cam_loc660[14:0]) |
 (snoop_in == cam_loc661[14:0]) |
 (snoop_in == cam_loc662[14:0]) |
 (snoop_in == cam_loc663[14:0]) |
 (snoop_in == cam_loc664[14:0]) |
 (snoop_in == cam_loc665[14:0]) |
 (snoop_in == cam_loc666[14:0]) |
 (snoop_in == cam_loc667[14:0]) |
 (snoop_in == cam_loc668[14:0]) |
 (snoop_in == cam_loc669[14:0]) |
 (snoop_in == cam_loc670[14:0]) |
 (snoop_in == cam_loc671[14:0]) |
 (snoop_in == cam_loc672[14:0]) |
 (snoop_in == cam_loc673[14:0]) |
 (snoop_in == cam_loc674[14:0]) |
 (snoop_in == cam_loc675[14:0]) |
 (snoop_in == cam_loc676[14:0]) |
 (snoop_in == cam_loc677[14:0]) |
 (snoop_in == cam_loc678[14:0]) |
 (snoop_in == cam_loc679[14:0]) |
 (snoop_in == cam_loc680[14:0]) |
 (snoop_in == cam_loc681[14:0]) |
 (snoop_in == cam_loc682[14:0]) |
 (snoop_in == cam_loc683[14:0]) |
 (snoop_in == cam_loc684[14:0]) |
 (snoop_in == cam_loc685[14:0]) |
 (snoop_in == cam_loc686[14:0]) |
 (snoop_in == cam_loc687[14:0]) |
 (snoop_in == cam_loc688[14:0]) |
 (snoop_in == cam_loc689[14:0]) |
 (snoop_in == cam_loc690[14:0]) |
 (snoop_in == cam_loc691[14:0]) |
 (snoop_in == cam_loc692[14:0]) |
 (snoop_in == cam_loc693[14:0]) |
 (snoop_in == cam_loc694[14:0]) |
 (snoop_in == cam_loc695[14:0]) |
 (snoop_in == cam_loc696[14:0]) |
 (snoop_in == cam_loc697[14:0]) |
 (snoop_in == cam_loc698[14:0]) |
 (snoop_in == cam_loc699[14:0]) |
 (snoop_in == cam_loc700[14:0]) |
 (snoop_in == cam_loc701[14:0]) |
 (snoop_in == cam_loc702[14:0]) |
 (snoop_in == cam_loc703[14:0]) |
 (snoop_in == cam_loc704[14:0]) |
 (snoop_in == cam_loc705[14:0]) |
 (snoop_in == cam_loc706[14:0]) |
 (snoop_in == cam_loc707[14:0]) |
 (snoop_in == cam_loc708[14:0]) |
 (snoop_in == cam_loc709[14:0]) |
 (snoop_in == cam_loc710[14:0]) |
 (snoop_in == cam_loc711[14:0]) |
 (snoop_in == cam_loc712[14:0]) |
 (snoop_in == cam_loc713[14:0]) |
 (snoop_in == cam_loc714[14:0]) |
 (snoop_in == cam_loc715[14:0]) |
 (snoop_in == cam_loc716[14:0]) |
 (snoop_in == cam_loc717[14:0]) |
 (snoop_in == cam_loc718[14:0]) |
 (snoop_in == cam_loc719[14:0]) |
 (snoop_in == cam_loc720[14:0]) |
 (snoop_in == cam_loc721[14:0]) |
 (snoop_in == cam_loc722[14:0]) |
 (snoop_in == cam_loc723[14:0]) |
 (snoop_in == cam_loc724[14:0]) |
 (snoop_in == cam_loc725[14:0]) |
 (snoop_in == cam_loc726[14:0]) |
 (snoop_in == cam_loc727[14:0]) |
 (snoop_in == cam_loc728[14:0]) |
 (snoop_in == cam_loc729[14:0]) |
 (snoop_in == cam_loc730[14:0]) |
 (snoop_in == cam_loc731[14:0]) |
 (snoop_in == cam_loc732[14:0]) |
 (snoop_in == cam_loc733[14:0]) |
 (snoop_in == cam_loc734[14:0]) |
 (snoop_in == cam_loc735[14:0]) |
 (snoop_in == cam_loc736[14:0]) |
 (snoop_in == cam_loc737[14:0]) |
 (snoop_in == cam_loc738[14:0]) |
 (snoop_in == cam_loc739[14:0]) |
 (snoop_in == cam_loc740[14:0]) |
 (snoop_in == cam_loc741[14:0]) |
 (snoop_in == cam_loc742[14:0]) |
 (snoop_in == cam_loc743[14:0]) |
 (snoop_in == cam_loc744[14:0]) |
 (snoop_in == cam_loc745[14:0]) |
 (snoop_in == cam_loc746[14:0]) |
 (snoop_in == cam_loc747[14:0]) |
 (snoop_in == cam_loc748[14:0]) |
 (snoop_in == cam_loc749[14:0]) |
 (snoop_in == cam_loc750[14:0]) |
 (snoop_in == cam_loc751[14:0]) |
 (snoop_in == cam_loc752[14:0]) |
 (snoop_in == cam_loc753[14:0]) |
 (snoop_in == cam_loc754[14:0]) |
 (snoop_in == cam_loc755[14:0]) |
 (snoop_in == cam_loc756[14:0]) |
 (snoop_in == cam_loc757[14:0]) |
 (snoop_in == cam_loc758[14:0]) |
 (snoop_in == cam_loc759[14:0]) |
 (snoop_in == cam_loc760[14:0]) |
 (snoop_in == cam_loc761[14:0]) |
 (snoop_in == cam_loc762[14:0]) |
 (snoop_in == cam_loc763[14:0]) |
 (snoop_in == cam_loc764[14:0]) |
 (snoop_in == cam_loc765[14:0]) |
 (snoop_in == cam_loc766[14:0]) |
 (snoop_in == cam_loc767[14:0]) |
 (snoop_in == cam_loc768[14:0]) |
 (snoop_in == cam_loc769[14:0]) |
 (snoop_in == cam_loc770[14:0]) |
 (snoop_in == cam_loc771[14:0]) |
 (snoop_in == cam_loc772[14:0]) |
 (snoop_in == cam_loc773[14:0]) |
 (snoop_in == cam_loc774[14:0]) |
 (snoop_in == cam_loc775[14:0]) |
 (snoop_in == cam_loc776[14:0]) |
 (snoop_in == cam_loc777[14:0]) |
 (snoop_in == cam_loc778[14:0]) |
 (snoop_in == cam_loc779[14:0]) |
 (snoop_in == cam_loc780[14:0]) |
 (snoop_in == cam_loc781[14:0]) |
 (snoop_in == cam_loc782[14:0]) |
 (snoop_in == cam_loc783[14:0]) |
 (snoop_in == cam_loc784[14:0]) |
 (snoop_in == cam_loc785[14:0]) |
 (snoop_in == cam_loc786[14:0]) |
 (snoop_in == cam_loc787[14:0]) |
 (snoop_in == cam_loc788[14:0]) |
 (snoop_in == cam_loc789[14:0]) |
 (snoop_in == cam_loc790[14:0]) |
 (snoop_in == cam_loc791[14:0]) |
 (snoop_in == cam_loc792[14:0]) |
 (snoop_in == cam_loc793[14:0]) |
 (snoop_in == cam_loc794[14:0]) |
 (snoop_in == cam_loc795[14:0]) |
 (snoop_in == cam_loc796[14:0]) |
 (snoop_in == cam_loc797[14:0]) |
 (snoop_in == cam_loc798[14:0]) |
 (snoop_in == cam_loc799[14:0]) |
 (snoop_in == cam_loc800[14:0]) |
 (snoop_in == cam_loc801[14:0]) |
 (snoop_in == cam_loc802[14:0]) |
 (snoop_in == cam_loc803[14:0]) |
 (snoop_in == cam_loc804[14:0]) |
 (snoop_in == cam_loc805[14:0]) |
 (snoop_in == cam_loc806[14:0]) |
 (snoop_in == cam_loc807[14:0]) |
 (snoop_in == cam_loc808[14:0]) |
 (snoop_in == cam_loc809[14:0]) |
 (snoop_in == cam_loc810[14:0]) |
 (snoop_in == cam_loc811[14:0]) |
 (snoop_in == cam_loc812[14:0]) |
 (snoop_in == cam_loc813[14:0]) |
 (snoop_in == cam_loc814[14:0]) |
 (snoop_in == cam_loc815[14:0]) |
 (snoop_in == cam_loc816[14:0]) |
 (snoop_in == cam_loc817[14:0]) |
 (snoop_in == cam_loc818[14:0]) |
 (snoop_in == cam_loc819[14:0]) |
 (snoop_in == cam_loc820[14:0]) |
 (snoop_in == cam_loc821[14:0]) |
 (snoop_in == cam_loc822[14:0]) |
 (snoop_in == cam_loc823[14:0]) |
 (snoop_in == cam_loc824[14:0]) |
 (snoop_in == cam_loc825[14:0]) |
 (snoop_in == cam_loc826[14:0]) |
 (snoop_in == cam_loc827[14:0]) |
 (snoop_in == cam_loc828[14:0]) |
 (snoop_in == cam_loc829[14:0]) |
 (snoop_in == cam_loc830[14:0]) |
 (snoop_in == cam_loc831[14:0]) |
 (snoop_in == cam_loc832[14:0]) |
 (snoop_in == cam_loc833[14:0]) |
 (snoop_in == cam_loc834[14:0]) |
 (snoop_in == cam_loc835[14:0]) |
 (snoop_in == cam_loc836[14:0]) |
 (snoop_in == cam_loc837[14:0]) |
 (snoop_in == cam_loc838[14:0]) |
 (snoop_in == cam_loc839[14:0]) |
 (snoop_in == cam_loc840[14:0]) |
 (snoop_in == cam_loc841[14:0]) |
 (snoop_in == cam_loc842[14:0]) |
 (snoop_in == cam_loc843[14:0]) |
 (snoop_in == cam_loc844[14:0]) |
 (snoop_in == cam_loc845[14:0]) |
 (snoop_in == cam_loc846[14:0]) |
 (snoop_in == cam_loc847[14:0]) |
 (snoop_in == cam_loc848[14:0]) |
 (snoop_in == cam_loc849[14:0]) |
 (snoop_in == cam_loc850[14:0]) |
 (snoop_in == cam_loc851[14:0]) |
 (snoop_in == cam_loc852[14:0]) |
 (snoop_in == cam_loc853[14:0]) |
 (snoop_in == cam_loc854[14:0]) |
 (snoop_in == cam_loc855[14:0]) |
 (snoop_in == cam_loc856[14:0]) |
 (snoop_in == cam_loc857[14:0]) |
 (snoop_in == cam_loc858[14:0]) |
 (snoop_in == cam_loc859[14:0]) |
 (snoop_in == cam_loc860[14:0]) |
 (snoop_in == cam_loc861[14:0]) |
 (snoop_in == cam_loc862[14:0]) |
 (snoop_in == cam_loc863[14:0]) |
 (snoop_in == cam_loc864[14:0]) |
 (snoop_in == cam_loc865[14:0]) |
 (snoop_in == cam_loc866[14:0]) |
 (snoop_in == cam_loc867[14:0]) |
 (snoop_in == cam_loc868[14:0]) |
 (snoop_in == cam_loc869[14:0]) |
 (snoop_in == cam_loc870[14:0]) |
 (snoop_in == cam_loc871[14:0]) |
 (snoop_in == cam_loc872[14:0]) |
 (snoop_in == cam_loc873[14:0]) |
 (snoop_in == cam_loc874[14:0]) |
 (snoop_in == cam_loc875[14:0]) |
 (snoop_in == cam_loc876[14:0]) |
 (snoop_in == cam_loc877[14:0]) |
 (snoop_in == cam_loc878[14:0]) |
 (snoop_in == cam_loc879[14:0]) |
 (snoop_in == cam_loc880[14:0]) |
 (snoop_in == cam_loc881[14:0]) |
 (snoop_in == cam_loc882[14:0]) |
 (snoop_in == cam_loc883[14:0]) |
 (snoop_in == cam_loc884[14:0]) |
 (snoop_in == cam_loc885[14:0]) |
 (snoop_in == cam_loc886[14:0]) |
 (snoop_in == cam_loc887[14:0]) |
 (snoop_in == cam_loc888[14:0]) |
 (snoop_in == cam_loc889[14:0]) |
 (snoop_in == cam_loc890[14:0]) |
 (snoop_in == cam_loc891[14:0]) |
 (snoop_in == cam_loc892[14:0]) |
 (snoop_in == cam_loc893[14:0]) |
 (snoop_in == cam_loc894[14:0]) |
 (snoop_in == cam_loc895[14:0]) |
 (snoop_in == cam_loc896[14:0]) |
 (snoop_in == cam_loc897[14:0]) |
 (snoop_in == cam_loc898[14:0]) |
 (snoop_in == cam_loc899[14:0]) |
 (snoop_in == cam_loc900[14:0]) |
 (snoop_in == cam_loc901[14:0]) |
 (snoop_in == cam_loc902[14:0]) |
 (snoop_in == cam_loc903[14:0]) |
 (snoop_in == cam_loc904[14:0]) |
 (snoop_in == cam_loc905[14:0]) |
 (snoop_in == cam_loc906[14:0]) |
 (snoop_in == cam_loc907[14:0]) |
 (snoop_in == cam_loc908[14:0]) |
 (snoop_in == cam_loc909[14:0]) |
 (snoop_in == cam_loc910[14:0]) |
 (snoop_in == cam_loc911[14:0]) |
 (snoop_in == cam_loc912[14:0]) |
 (snoop_in == cam_loc913[14:0]) |
 (snoop_in == cam_loc914[14:0]) |
 (snoop_in == cam_loc915[14:0]) |
 (snoop_in == cam_loc916[14:0]) |
 (snoop_in == cam_loc917[14:0]) |
 (snoop_in == cam_loc918[14:0]) |
 (snoop_in == cam_loc919[14:0]) |
 (snoop_in == cam_loc920[14:0]) |
 (snoop_in == cam_loc921[14:0]) |
 (snoop_in == cam_loc922[14:0]) |
 (snoop_in == cam_loc923[14:0]) |
 (snoop_in == cam_loc924[14:0]) |
 (snoop_in == cam_loc925[14:0]) |
 (snoop_in == cam_loc926[14:0]) |
 (snoop_in == cam_loc927[14:0]) |
 (snoop_in == cam_loc928[14:0]) |
 (snoop_in == cam_loc929[14:0]) |
 (snoop_in == cam_loc930[14:0]) |
 (snoop_in == cam_loc931[14:0]) |
 (snoop_in == cam_loc932[14:0]) |
 (snoop_in == cam_loc933[14:0]) |
 (snoop_in == cam_loc934[14:0]) |
 (snoop_in == cam_loc935[14:0]) |
 (snoop_in == cam_loc936[14:0]) |
 (snoop_in == cam_loc937[14:0]) |
 (snoop_in == cam_loc938[14:0]) |
 (snoop_in == cam_loc939[14:0]) |
 (snoop_in == cam_loc940[14:0]) |
 (snoop_in == cam_loc941[14:0]) |
 (snoop_in == cam_loc942[14:0]) |
 (snoop_in == cam_loc943[14:0]) |
 (snoop_in == cam_loc944[14:0]) |
 (snoop_in == cam_loc945[14:0]) |
 (snoop_in == cam_loc946[14:0]) |
 (snoop_in == cam_loc947[14:0]) |
 (snoop_in == cam_loc948[14:0]) |
 (snoop_in == cam_loc949[14:0]) |
 (snoop_in == cam_loc950[14:0]) |
 (snoop_in == cam_loc951[14:0]) |
 (snoop_in == cam_loc952[14:0]) |
 (snoop_in == cam_loc953[14:0]) |
 (snoop_in == cam_loc954[14:0]) |
 (snoop_in == cam_loc955[14:0]) |
 (snoop_in == cam_loc956[14:0]) |
 (snoop_in == cam_loc957[14:0]) |
 (snoop_in == cam_loc958[14:0]) |
 (snoop_in == cam_loc959[14:0]) |
 (snoop_in == cam_loc960[14:0]) |
 (snoop_in == cam_loc961[14:0]) |
 (snoop_in == cam_loc962[14:0]) |
 (snoop_in == cam_loc963[14:0]) |
 (snoop_in == cam_loc964[14:0]) |
 (snoop_in == cam_loc965[14:0]) |
 (snoop_in == cam_loc966[14:0]) |
 (snoop_in == cam_loc967[14:0]) |
 (snoop_in == cam_loc968[14:0]) |
 (snoop_in == cam_loc969[14:0]) |
 (snoop_in == cam_loc970[14:0]) |
 (snoop_in == cam_loc971[14:0]) |
 (snoop_in == cam_loc972[14:0]) |
 (snoop_in == cam_loc973[14:0]) |
 (snoop_in == cam_loc974[14:0]) |
 (snoop_in == cam_loc975[14:0]) |
 (snoop_in == cam_loc976[14:0]) |
 (snoop_in == cam_loc977[14:0]) |
 (snoop_in == cam_loc978[14:0]) |
 (snoop_in == cam_loc979[14:0]) |
 (snoop_in == cam_loc980[14:0]) |
 (snoop_in == cam_loc981[14:0]) |
 (snoop_in == cam_loc982[14:0]) |
 (snoop_in == cam_loc983[14:0]) |
 (snoop_in == cam_loc984[14:0]) |
 (snoop_in == cam_loc985[14:0]) |
 (snoop_in == cam_loc986[14:0]) |
 (snoop_in == cam_loc987[14:0]) |
 (snoop_in == cam_loc988[14:0]) |
 (snoop_in == cam_loc989[14:0]) |
 (snoop_in == cam_loc990[14:0]) |
 (snoop_in == cam_loc991[14:0]) |
 (snoop_in == cam_loc992[14:0]) |
 (snoop_in == cam_loc993[14:0]) |
 (snoop_in == cam_loc994[14:0]) |
 (snoop_in == cam_loc995[14:0]) |
 (snoop_in == cam_loc996[14:0]) |
 (snoop_in == cam_loc997[14:0]) |
 (snoop_in == cam_loc998[14:0]) |
 (snoop_in == cam_loc999[14:0]) |
 (snoop_in == cam_loc1000[14:0]) |
 (snoop_in == cam_loc1001[14:0]) |
 (snoop_in == cam_loc1002[14:0]) |
 (snoop_in == cam_loc1003[14:0]) |
 (snoop_in == cam_loc1004[14:0]) |
 (snoop_in == cam_loc1005[14:0]) |
 (snoop_in == cam_loc1006[14:0]) |
 (snoop_in == cam_loc1007[14:0]) |
 (snoop_in == cam_loc1008[14:0]) |
 (snoop_in == cam_loc1009[14:0]) |
 (snoop_in == cam_loc1010[14:0]) |
 (snoop_in == cam_loc1011[14:0]) |
 (snoop_in == cam_loc1012[14:0]) |
 (snoop_in == cam_loc1013[14:0]) |
 (snoop_in == cam_loc1014[14:0]) |
 (snoop_in == cam_loc1015[14:0]) |
 (snoop_in == cam_loc1016[14:0]) |
 (snoop_in == cam_loc1017[14:0]) |
 (snoop_in == cam_loc1018[14:0]) |
 (snoop_in == cam_loc1019[14:0]) |
 (snoop_in == cam_loc1020[14:0]) |
 (snoop_in == cam_loc1021[14:0]) |
 (snoop_in == cam_loc1022[14:0]) |
 (snoop_in == cam_loc1023[14:0]) |
 (snoop_in == cam_loc1024[14:0]) |
 (snoop_in == cam_loc1025[14:0]) |
 (snoop_in == cam_loc1026[14:0]) |
 (snoop_in == cam_loc1027[14:0]) |
 (snoop_in == cam_loc1028[14:0]) |
 (snoop_in == cam_loc1029[14:0]) |
 (snoop_in == cam_loc1030[14:0]) |
 (snoop_in == cam_loc1031[14:0]) |
 (snoop_in == cam_loc1032[14:0]) |
 (snoop_in == cam_loc1033[14:0]) |
 (snoop_in == cam_loc1034[14:0]) |
 (snoop_in == cam_loc1035[14:0]) |
 (snoop_in == cam_loc1036[14:0]) |
 (snoop_in == cam_loc1037[14:0]) |
 (snoop_in == cam_loc1038[14:0]) |
 (snoop_in == cam_loc1039[14:0]) |
 (snoop_in == cam_loc1040[14:0]) |
 (snoop_in == cam_loc1041[14:0]) |
 (snoop_in == cam_loc1042[14:0]) |
 (snoop_in == cam_loc1043[14:0]) |
 (snoop_in == cam_loc1044[14:0]) |
 (snoop_in == cam_loc1045[14:0]) |
 (snoop_in == cam_loc1046[14:0]) |
 (snoop_in == cam_loc1047[14:0]) |
 (snoop_in == cam_loc1048[14:0]) |
 (snoop_in == cam_loc1049[14:0]) |
 (snoop_in == cam_loc1050[14:0]) |
 (snoop_in == cam_loc1051[14:0]) |
 (snoop_in == cam_loc1052[14:0]) |
 (snoop_in == cam_loc1053[14:0]) |
 (snoop_in == cam_loc1054[14:0]) |
 (snoop_in == cam_loc1055[14:0]) |
 (snoop_in == cam_loc1056[14:0]) |
 (snoop_in == cam_loc1057[14:0]) |
 (snoop_in == cam_loc1058[14:0]) |
 (snoop_in == cam_loc1059[14:0]) |
 (snoop_in == cam_loc1060[14:0]) |
 (snoop_in == cam_loc1061[14:0]) |
 (snoop_in == cam_loc1062[14:0]) |
 (snoop_in == cam_loc1063[14:0]) |
 (snoop_in == cam_loc1064[14:0]) |
 (snoop_in == cam_loc1065[14:0]) |
 (snoop_in == cam_loc1066[14:0]) |
 (snoop_in == cam_loc1067[14:0]) |
 (snoop_in == cam_loc1068[14:0]) |
 (snoop_in == cam_loc1069[14:0]) |
 (snoop_in == cam_loc1070[14:0]) |
 (snoop_in == cam_loc1071[14:0]) |
 (snoop_in == cam_loc1072[14:0]) |
 (snoop_in == cam_loc1073[14:0]) |
 (snoop_in == cam_loc1074[14:0]) |
 (snoop_in == cam_loc1075[14:0]) |
 (snoop_in == cam_loc1076[14:0]) |
 (snoop_in == cam_loc1077[14:0]) |
 (snoop_in == cam_loc1078[14:0]) |
 (snoop_in == cam_loc1079[14:0]) |
 (snoop_in == cam_loc1080[14:0]) |
 (snoop_in == cam_loc1081[14:0]) |
 (snoop_in == cam_loc1082[14:0]) |
 (snoop_in == cam_loc1083[14:0]) |
 (snoop_in == cam_loc1084[14:0]) |
 (snoop_in == cam_loc1085[14:0]) |
 (snoop_in == cam_loc1086[14:0]) |
 (snoop_in == cam_loc1087[14:0]) |
 (snoop_in == cam_loc1088[14:0]) |
 (snoop_in == cam_loc1089[14:0]) |
 (snoop_in == cam_loc1090[14:0]) |
 (snoop_in == cam_loc1091[14:0]) |
 (snoop_in == cam_loc1092[14:0]) |
 (snoop_in == cam_loc1093[14:0]) |
 (snoop_in == cam_loc1094[14:0]) |
 (snoop_in == cam_loc1095[14:0]) |
 (snoop_in == cam_loc1096[14:0]) |
 (snoop_in == cam_loc1097[14:0]) |
 (snoop_in == cam_loc1098[14:0]) |
 (snoop_in == cam_loc1099[14:0])

);

wire assign snoop_data = 20'd0 |
( (snoop_in == cam_loc0[14:0]) ? cam_loc0 : 20'd0 ) |
 ( (snoop_in == cam_loc1[14:0]) ? cam_loc1 : 20'd0 ) |
 ( (snoop_in == cam_loc2[14:0]) ? cam_loc2 : 20'd0 ) |
 ( (snoop_in == cam_loc3[14:0]) ? cam_loc3 : 20'd0 ) |
 ( (snoop_in == cam_loc4[14:0]) ? cam_loc4 : 20'd0 ) |
 ( (snoop_in == cam_loc5[14:0]) ? cam_loc5 : 20'd0 ) |
 ( (snoop_in == cam_loc6[14:0]) ? cam_loc6 : 20'd0 ) |
 ( (snoop_in == cam_loc7[14:0]) ? cam_loc7 : 20'd0 ) |
 ( (snoop_in == cam_loc8[14:0]) ? cam_loc8 : 20'd0 ) |
 ( (snoop_in == cam_loc9[14:0]) ? cam_loc9 : 20'd0 ) |
 ( (snoop_in == cam_loc10[14:0]) ? cam_loc10 : 20'd0 ) |
 ( (snoop_in == cam_loc11[14:0]) ? cam_loc11 : 20'd0 ) |
 ( (snoop_in == cam_loc12[14:0]) ? cam_loc12 : 20'd0 ) |
 ( (snoop_in == cam_loc13[14:0]) ? cam_loc13 : 20'd0 ) |
 ( (snoop_in == cam_loc14[14:0]) ? cam_loc14 : 20'd0 ) |
 ( (snoop_in == cam_loc15[14:0]) ? cam_loc15 : 20'd0 ) |
 ( (snoop_in == cam_loc16[14:0]) ? cam_loc16 : 20'd0 ) |
 ( (snoop_in == cam_loc17[14:0]) ? cam_loc17 : 20'd0 ) |
 ( (snoop_in == cam_loc18[14:0]) ? cam_loc18 : 20'd0 ) |
 ( (snoop_in == cam_loc19[14:0]) ? cam_loc19 : 20'd0 ) |
 ( (snoop_in == cam_loc20[14:0]) ? cam_loc20 : 20'd0 ) |
 ( (snoop_in == cam_loc21[14:0]) ? cam_loc21 : 20'd0 ) |
 ( (snoop_in == cam_loc22[14:0]) ? cam_loc22 : 20'd0 ) |
 ( (snoop_in == cam_loc23[14:0]) ? cam_loc23 : 20'd0 ) |
 ( (snoop_in == cam_loc24[14:0]) ? cam_loc24 : 20'd0 ) |
 ( (snoop_in == cam_loc25[14:0]) ? cam_loc25 : 20'd0 ) |
 ( (snoop_in == cam_loc26[14:0]) ? cam_loc26 : 20'd0 ) |
 ( (snoop_in == cam_loc27[14:0]) ? cam_loc27 : 20'd0 ) |
 ( (snoop_in == cam_loc28[14:0]) ? cam_loc28 : 20'd0 ) |
 ( (snoop_in == cam_loc29[14:0]) ? cam_loc29 : 20'd0 ) |
 ( (snoop_in == cam_loc30[14:0]) ? cam_loc30 : 20'd0 ) |
 ( (snoop_in == cam_loc31[14:0]) ? cam_loc31 : 20'd0 ) |
 ( (snoop_in == cam_loc32[14:0]) ? cam_loc32 : 20'd0 ) |
 ( (snoop_in == cam_loc33[14:0]) ? cam_loc33 : 20'd0 ) |
 ( (snoop_in == cam_loc34[14:0]) ? cam_loc34 : 20'd0 ) |
 ( (snoop_in == cam_loc35[14:0]) ? cam_loc35 : 20'd0 ) |
 ( (snoop_in == cam_loc36[14:0]) ? cam_loc36 : 20'd0 ) |
 ( (snoop_in == cam_loc37[14:0]) ? cam_loc37 : 20'd0 ) |
 ( (snoop_in == cam_loc38[14:0]) ? cam_loc38 : 20'd0 ) |
 ( (snoop_in == cam_loc39[14:0]) ? cam_loc39 : 20'd0 ) |
 ( (snoop_in == cam_loc40[14:0]) ? cam_loc40 : 20'd0 ) |
 ( (snoop_in == cam_loc41[14:0]) ? cam_loc41 : 20'd0 ) |
 ( (snoop_in == cam_loc42[14:0]) ? cam_loc42 : 20'd0 ) |
 ( (snoop_in == cam_loc43[14:0]) ? cam_loc43 : 20'd0 ) |
 ( (snoop_in == cam_loc44[14:0]) ? cam_loc44 : 20'd0 ) |
 ( (snoop_in == cam_loc45[14:0]) ? cam_loc45 : 20'd0 ) |
 ( (snoop_in == cam_loc46[14:0]) ? cam_loc46 : 20'd0 ) |
 ( (snoop_in == cam_loc47[14:0]) ? cam_loc47 : 20'd0 ) |
 ( (snoop_in == cam_loc48[14:0]) ? cam_loc48 : 20'd0 ) |
 ( (snoop_in == cam_loc49[14:0]) ? cam_loc49 : 20'd0 ) |
 ( (snoop_in == cam_loc50[14:0]) ? cam_loc50 : 20'd0 ) |
 ( (snoop_in == cam_loc51[14:0]) ? cam_loc51 : 20'd0 ) |
 ( (snoop_in == cam_loc52[14:0]) ? cam_loc52 : 20'd0 ) |
 ( (snoop_in == cam_loc53[14:0]) ? cam_loc53 : 20'd0 ) |
 ( (snoop_in == cam_loc54[14:0]) ? cam_loc54 : 20'd0 ) |
 ( (snoop_in == cam_loc55[14:0]) ? cam_loc55 : 20'd0 ) |
 ( (snoop_in == cam_loc56[14:0]) ? cam_loc56 : 20'd0 ) |
 ( (snoop_in == cam_loc57[14:0]) ? cam_loc57 : 20'd0 ) |
 ( (snoop_in == cam_loc58[14:0]) ? cam_loc58 : 20'd0 ) |
 ( (snoop_in == cam_loc59[14:0]) ? cam_loc59 : 20'd0 ) |
 ( (snoop_in == cam_loc60[14:0]) ? cam_loc60 : 20'd0 ) |
 ( (snoop_in == cam_loc61[14:0]) ? cam_loc61 : 20'd0 ) |
 ( (snoop_in == cam_loc62[14:0]) ? cam_loc62 : 20'd0 ) |
 ( (snoop_in == cam_loc63[14:0]) ? cam_loc63 : 20'd0 ) |
 ( (snoop_in == cam_loc64[14:0]) ? cam_loc64 : 20'd0 ) |
 ( (snoop_in == cam_loc65[14:0]) ? cam_loc65 : 20'd0 ) |
 ( (snoop_in == cam_loc66[14:0]) ? cam_loc66 : 20'd0 ) |
 ( (snoop_in == cam_loc67[14:0]) ? cam_loc67 : 20'd0 ) |
 ( (snoop_in == cam_loc68[14:0]) ? cam_loc68 : 20'd0 ) |
 ( (snoop_in == cam_loc69[14:0]) ? cam_loc69 : 20'd0 ) |
 ( (snoop_in == cam_loc70[14:0]) ? cam_loc70 : 20'd0 ) |
 ( (snoop_in == cam_loc71[14:0]) ? cam_loc71 : 20'd0 ) |
 ( (snoop_in == cam_loc72[14:0]) ? cam_loc72 : 20'd0 ) |
 ( (snoop_in == cam_loc73[14:0]) ? cam_loc73 : 20'd0 ) |
 ( (snoop_in == cam_loc74[14:0]) ? cam_loc74 : 20'd0 ) |
 ( (snoop_in == cam_loc75[14:0]) ? cam_loc75 : 20'd0 ) |
 ( (snoop_in == cam_loc76[14:0]) ? cam_loc76 : 20'd0 ) |
 ( (snoop_in == cam_loc77[14:0]) ? cam_loc77 : 20'd0 ) |
 ( (snoop_in == cam_loc78[14:0]) ? cam_loc78 : 20'd0 ) |
 ( (snoop_in == cam_loc79[14:0]) ? cam_loc79 : 20'd0 ) |
 ( (snoop_in == cam_loc80[14:0]) ? cam_loc80 : 20'd0 ) |
 ( (snoop_in == cam_loc81[14:0]) ? cam_loc81 : 20'd0 ) |
 ( (snoop_in == cam_loc82[14:0]) ? cam_loc82 : 20'd0 ) |
 ( (snoop_in == cam_loc83[14:0]) ? cam_loc83 : 20'd0 ) |
 ( (snoop_in == cam_loc84[14:0]) ? cam_loc84 : 20'd0 ) |
 ( (snoop_in == cam_loc85[14:0]) ? cam_loc85 : 20'd0 ) |
 ( (snoop_in == cam_loc86[14:0]) ? cam_loc86 : 20'd0 ) |
 ( (snoop_in == cam_loc87[14:0]) ? cam_loc87 : 20'd0 ) |
 ( (snoop_in == cam_loc88[14:0]) ? cam_loc88 : 20'd0 ) |
 ( (snoop_in == cam_loc89[14:0]) ? cam_loc89 : 20'd0 ) |
 ( (snoop_in == cam_loc90[14:0]) ? cam_loc90 : 20'd0 ) |
 ( (snoop_in == cam_loc91[14:0]) ? cam_loc91 : 20'd0 ) |
 ( (snoop_in == cam_loc92[14:0]) ? cam_loc92 : 20'd0 ) |
 ( (snoop_in == cam_loc93[14:0]) ? cam_loc93 : 20'd0 ) |
 ( (snoop_in == cam_loc94[14:0]) ? cam_loc94 : 20'd0 ) |
 ( (snoop_in == cam_loc95[14:0]) ? cam_loc95 : 20'd0 ) |
 ( (snoop_in == cam_loc96[14:0]) ? cam_loc96 : 20'd0 ) |
 ( (snoop_in == cam_loc97[14:0]) ? cam_loc97 : 20'd0 ) |
 ( (snoop_in == cam_loc98[14:0]) ? cam_loc98 : 20'd0 ) |
 ( (snoop_in == cam_loc99[14:0]) ? cam_loc99 : 20'd0 ) |
 ( (snoop_in == cam_loc100[14:0]) ? cam_loc100 : 20'd0 ) |
 ( (snoop_in == cam_loc101[14:0]) ? cam_loc101 : 20'd0 ) |
 ( (snoop_in == cam_loc102[14:0]) ? cam_loc102 : 20'd0 ) |
 ( (snoop_in == cam_loc103[14:0]) ? cam_loc103 : 20'd0 ) |
 ( (snoop_in == cam_loc104[14:0]) ? cam_loc104 : 20'd0 ) |
 ( (snoop_in == cam_loc105[14:0]) ? cam_loc105 : 20'd0 ) |
 ( (snoop_in == cam_loc106[14:0]) ? cam_loc106 : 20'd0 ) |
 ( (snoop_in == cam_loc107[14:0]) ? cam_loc107 : 20'd0 ) |
 ( (snoop_in == cam_loc108[14:0]) ? cam_loc108 : 20'd0 ) |
 ( (snoop_in == cam_loc109[14:0]) ? cam_loc109 : 20'd0 ) |
 ( (snoop_in == cam_loc110[14:0]) ? cam_loc110 : 20'd0 ) |
 ( (snoop_in == cam_loc111[14:0]) ? cam_loc111 : 20'd0 ) |
 ( (snoop_in == cam_loc112[14:0]) ? cam_loc112 : 20'd0 ) |
 ( (snoop_in == cam_loc113[14:0]) ? cam_loc113 : 20'd0 ) |
 ( (snoop_in == cam_loc114[14:0]) ? cam_loc114 : 20'd0 ) |
 ( (snoop_in == cam_loc115[14:0]) ? cam_loc115 : 20'd0 ) |
 ( (snoop_in == cam_loc116[14:0]) ? cam_loc116 : 20'd0 ) |
 ( (snoop_in == cam_loc117[14:0]) ? cam_loc117 : 20'd0 ) |
 ( (snoop_in == cam_loc118[14:0]) ? cam_loc118 : 20'd0 ) |
 ( (snoop_in == cam_loc119[14:0]) ? cam_loc119 : 20'd0 ) |
 ( (snoop_in == cam_loc120[14:0]) ? cam_loc120 : 20'd0 ) |
 ( (snoop_in == cam_loc121[14:0]) ? cam_loc121 : 20'd0 ) |
 ( (snoop_in == cam_loc122[14:0]) ? cam_loc122 : 20'd0 ) |
 ( (snoop_in == cam_loc123[14:0]) ? cam_loc123 : 20'd0 ) |
 ( (snoop_in == cam_loc124[14:0]) ? cam_loc124 : 20'd0 ) |
 ( (snoop_in == cam_loc125[14:0]) ? cam_loc125 : 20'd0 ) |
 ( (snoop_in == cam_loc126[14:0]) ? cam_loc126 : 20'd0 ) |
 ( (snoop_in == cam_loc127[14:0]) ? cam_loc127 : 20'd0 ) |
 ( (snoop_in == cam_loc128[14:0]) ? cam_loc128 : 20'd0 ) |
 ( (snoop_in == cam_loc129[14:0]) ? cam_loc129 : 20'd0 ) |
 ( (snoop_in == cam_loc130[14:0]) ? cam_loc130 : 20'd0 ) |
 ( (snoop_in == cam_loc131[14:0]) ? cam_loc131 : 20'd0 ) |
 ( (snoop_in == cam_loc132[14:0]) ? cam_loc132 : 20'd0 ) |
 ( (snoop_in == cam_loc133[14:0]) ? cam_loc133 : 20'd0 ) |
 ( (snoop_in == cam_loc134[14:0]) ? cam_loc134 : 20'd0 ) |
 ( (snoop_in == cam_loc135[14:0]) ? cam_loc135 : 20'd0 ) |
 ( (snoop_in == cam_loc136[14:0]) ? cam_loc136 : 20'd0 ) |
 ( (snoop_in == cam_loc137[14:0]) ? cam_loc137 : 20'd0 ) |
 ( (snoop_in == cam_loc138[14:0]) ? cam_loc138 : 20'd0 ) |
 ( (snoop_in == cam_loc139[14:0]) ? cam_loc139 : 20'd0 ) |
 ( (snoop_in == cam_loc140[14:0]) ? cam_loc140 : 20'd0 ) |
 ( (snoop_in == cam_loc141[14:0]) ? cam_loc141 : 20'd0 ) |
 ( (snoop_in == cam_loc142[14:0]) ? cam_loc142 : 20'd0 ) |
 ( (snoop_in == cam_loc143[14:0]) ? cam_loc143 : 20'd0 ) |
 ( (snoop_in == cam_loc144[14:0]) ? cam_loc144 : 20'd0 ) |
 ( (snoop_in == cam_loc145[14:0]) ? cam_loc145 : 20'd0 ) |
 ( (snoop_in == cam_loc146[14:0]) ? cam_loc146 : 20'd0 ) |
 ( (snoop_in == cam_loc147[14:0]) ? cam_loc147 : 20'd0 ) |
 ( (snoop_in == cam_loc148[14:0]) ? cam_loc148 : 20'd0 ) |
 ( (snoop_in == cam_loc149[14:0]) ? cam_loc149 : 20'd0 ) |
 ( (snoop_in == cam_loc150[14:0]) ? cam_loc150 : 20'd0 ) |
 ( (snoop_in == cam_loc151[14:0]) ? cam_loc151 : 20'd0 ) |
 ( (snoop_in == cam_loc152[14:0]) ? cam_loc152 : 20'd0 ) |
 ( (snoop_in == cam_loc153[14:0]) ? cam_loc153 : 20'd0 ) |
 ( (snoop_in == cam_loc154[14:0]) ? cam_loc154 : 20'd0 ) |
 ( (snoop_in == cam_loc155[14:0]) ? cam_loc155 : 20'd0 ) |
 ( (snoop_in == cam_loc156[14:0]) ? cam_loc156 : 20'd0 ) |
 ( (snoop_in == cam_loc157[14:0]) ? cam_loc157 : 20'd0 ) |
 ( (snoop_in == cam_loc158[14:0]) ? cam_loc158 : 20'd0 ) |
 ( (snoop_in == cam_loc159[14:0]) ? cam_loc159 : 20'd0 ) |
 ( (snoop_in == cam_loc160[14:0]) ? cam_loc160 : 20'd0 ) |
 ( (snoop_in == cam_loc161[14:0]) ? cam_loc161 : 20'd0 ) |
 ( (snoop_in == cam_loc162[14:0]) ? cam_loc162 : 20'd0 ) |
 ( (snoop_in == cam_loc163[14:0]) ? cam_loc163 : 20'd0 ) |
 ( (snoop_in == cam_loc164[14:0]) ? cam_loc164 : 20'd0 ) |
 ( (snoop_in == cam_loc165[14:0]) ? cam_loc165 : 20'd0 ) |
 ( (snoop_in == cam_loc166[14:0]) ? cam_loc166 : 20'd0 ) |
 ( (snoop_in == cam_loc167[14:0]) ? cam_loc167 : 20'd0 ) |
 ( (snoop_in == cam_loc168[14:0]) ? cam_loc168 : 20'd0 ) |
 ( (snoop_in == cam_loc169[14:0]) ? cam_loc169 : 20'd0 ) |
 ( (snoop_in == cam_loc170[14:0]) ? cam_loc170 : 20'd0 ) |
 ( (snoop_in == cam_loc171[14:0]) ? cam_loc171 : 20'd0 ) |
 ( (snoop_in == cam_loc172[14:0]) ? cam_loc172 : 20'd0 ) |
 ( (snoop_in == cam_loc173[14:0]) ? cam_loc173 : 20'd0 ) |
 ( (snoop_in == cam_loc174[14:0]) ? cam_loc174 : 20'd0 ) |
 ( (snoop_in == cam_loc175[14:0]) ? cam_loc175 : 20'd0 ) |
 ( (snoop_in == cam_loc176[14:0]) ? cam_loc176 : 20'd0 ) |
 ( (snoop_in == cam_loc177[14:0]) ? cam_loc177 : 20'd0 ) |
 ( (snoop_in == cam_loc178[14:0]) ? cam_loc178 : 20'd0 ) |
 ( (snoop_in == cam_loc179[14:0]) ? cam_loc179 : 20'd0 ) |
 ( (snoop_in == cam_loc180[14:0]) ? cam_loc180 : 20'd0 ) |
 ( (snoop_in == cam_loc181[14:0]) ? cam_loc181 : 20'd0 ) |
 ( (snoop_in == cam_loc182[14:0]) ? cam_loc182 : 20'd0 ) |
 ( (snoop_in == cam_loc183[14:0]) ? cam_loc183 : 20'd0 ) |
 ( (snoop_in == cam_loc184[14:0]) ? cam_loc184 : 20'd0 ) |
 ( (snoop_in == cam_loc185[14:0]) ? cam_loc185 : 20'd0 ) |
 ( (snoop_in == cam_loc186[14:0]) ? cam_loc186 : 20'd0 ) |
 ( (snoop_in == cam_loc187[14:0]) ? cam_loc187 : 20'd0 ) |
 ( (snoop_in == cam_loc188[14:0]) ? cam_loc188 : 20'd0 ) |
 ( (snoop_in == cam_loc189[14:0]) ? cam_loc189 : 20'd0 ) |
 ( (snoop_in == cam_loc190[14:0]) ? cam_loc190 : 20'd0 ) |
 ( (snoop_in == cam_loc191[14:0]) ? cam_loc191 : 20'd0 ) |
 ( (snoop_in == cam_loc192[14:0]) ? cam_loc192 : 20'd0 ) |
 ( (snoop_in == cam_loc193[14:0]) ? cam_loc193 : 20'd0 ) |
 ( (snoop_in == cam_loc194[14:0]) ? cam_loc194 : 20'd0 ) |
 ( (snoop_in == cam_loc195[14:0]) ? cam_loc195 : 20'd0 ) |
 ( (snoop_in == cam_loc196[14:0]) ? cam_loc196 : 20'd0 ) |
 ( (snoop_in == cam_loc197[14:0]) ? cam_loc197 : 20'd0 ) |
 ( (snoop_in == cam_loc198[14:0]) ? cam_loc198 : 20'd0 ) |
 ( (snoop_in == cam_loc199[14:0]) ? cam_loc199 : 20'd0 ) |
 ( (snoop_in == cam_loc200[14:0]) ? cam_loc200 : 20'd0 ) |
 ( (snoop_in == cam_loc201[14:0]) ? cam_loc201 : 20'd0 ) |
 ( (snoop_in == cam_loc202[14:0]) ? cam_loc202 : 20'd0 ) |
 ( (snoop_in == cam_loc203[14:0]) ? cam_loc203 : 20'd0 ) |
 ( (snoop_in == cam_loc204[14:0]) ? cam_loc204 : 20'd0 ) |
 ( (snoop_in == cam_loc205[14:0]) ? cam_loc205 : 20'd0 ) |
 ( (snoop_in == cam_loc206[14:0]) ? cam_loc206 : 20'd0 ) |
 ( (snoop_in == cam_loc207[14:0]) ? cam_loc207 : 20'd0 ) |
 ( (snoop_in == cam_loc208[14:0]) ? cam_loc208 : 20'd0 ) |
 ( (snoop_in == cam_loc209[14:0]) ? cam_loc209 : 20'd0 ) |
 ( (snoop_in == cam_loc210[14:0]) ? cam_loc210 : 20'd0 ) |
 ( (snoop_in == cam_loc211[14:0]) ? cam_loc211 : 20'd0 ) |
 ( (snoop_in == cam_loc212[14:0]) ? cam_loc212 : 20'd0 ) |
 ( (snoop_in == cam_loc213[14:0]) ? cam_loc213 : 20'd0 ) |
 ( (snoop_in == cam_loc214[14:0]) ? cam_loc214 : 20'd0 ) |
 ( (snoop_in == cam_loc215[14:0]) ? cam_loc215 : 20'd0 ) |
 ( (snoop_in == cam_loc216[14:0]) ? cam_loc216 : 20'd0 ) |
 ( (snoop_in == cam_loc217[14:0]) ? cam_loc217 : 20'd0 ) |
 ( (snoop_in == cam_loc218[14:0]) ? cam_loc218 : 20'd0 ) |
 ( (snoop_in == cam_loc219[14:0]) ? cam_loc219 : 20'd0 ) |
 ( (snoop_in == cam_loc220[14:0]) ? cam_loc220 : 20'd0 ) |
 ( (snoop_in == cam_loc221[14:0]) ? cam_loc221 : 20'd0 ) |
 ( (snoop_in == cam_loc222[14:0]) ? cam_loc222 : 20'd0 ) |
 ( (snoop_in == cam_loc223[14:0]) ? cam_loc223 : 20'd0 ) |
 ( (snoop_in == cam_loc224[14:0]) ? cam_loc224 : 20'd0 ) |
 ( (snoop_in == cam_loc225[14:0]) ? cam_loc225 : 20'd0 ) |
 ( (snoop_in == cam_loc226[14:0]) ? cam_loc226 : 20'd0 ) |
 ( (snoop_in == cam_loc227[14:0]) ? cam_loc227 : 20'd0 ) |
 ( (snoop_in == cam_loc228[14:0]) ? cam_loc228 : 20'd0 ) |
 ( (snoop_in == cam_loc229[14:0]) ? cam_loc229 : 20'd0 ) |
 ( (snoop_in == cam_loc230[14:0]) ? cam_loc230 : 20'd0 ) |
 ( (snoop_in == cam_loc231[14:0]) ? cam_loc231 : 20'd0 ) |
 ( (snoop_in == cam_loc232[14:0]) ? cam_loc232 : 20'd0 ) |
 ( (snoop_in == cam_loc233[14:0]) ? cam_loc233 : 20'd0 ) |
 ( (snoop_in == cam_loc234[14:0]) ? cam_loc234 : 20'd0 ) |
 ( (snoop_in == cam_loc235[14:0]) ? cam_loc235 : 20'd0 ) |
 ( (snoop_in == cam_loc236[14:0]) ? cam_loc236 : 20'd0 ) |
 ( (snoop_in == cam_loc237[14:0]) ? cam_loc237 : 20'd0 ) |
 ( (snoop_in == cam_loc238[14:0]) ? cam_loc238 : 20'd0 ) |
 ( (snoop_in == cam_loc239[14:0]) ? cam_loc239 : 20'd0 ) |
 ( (snoop_in == cam_loc240[14:0]) ? cam_loc240 : 20'd0 ) |
 ( (snoop_in == cam_loc241[14:0]) ? cam_loc241 : 20'd0 ) |
 ( (snoop_in == cam_loc242[14:0]) ? cam_loc242 : 20'd0 ) |
 ( (snoop_in == cam_loc243[14:0]) ? cam_loc243 : 20'd0 ) |
 ( (snoop_in == cam_loc244[14:0]) ? cam_loc244 : 20'd0 ) |
 ( (snoop_in == cam_loc245[14:0]) ? cam_loc245 : 20'd0 ) |
 ( (snoop_in == cam_loc246[14:0]) ? cam_loc246 : 20'd0 ) |
 ( (snoop_in == cam_loc247[14:0]) ? cam_loc247 : 20'd0 ) |
 ( (snoop_in == cam_loc248[14:0]) ? cam_loc248 : 20'd0 ) |
 ( (snoop_in == cam_loc249[14:0]) ? cam_loc249 : 20'd0 ) |
 ( (snoop_in == cam_loc250[14:0]) ? cam_loc250 : 20'd0 ) |
 ( (snoop_in == cam_loc251[14:0]) ? cam_loc251 : 20'd0 ) |
 ( (snoop_in == cam_loc252[14:0]) ? cam_loc252 : 20'd0 ) |
 ( (snoop_in == cam_loc253[14:0]) ? cam_loc253 : 20'd0 ) |
 ( (snoop_in == cam_loc254[14:0]) ? cam_loc254 : 20'd0 ) |
 ( (snoop_in == cam_loc255[14:0]) ? cam_loc255 : 20'd0 ) |
 ( (snoop_in == cam_loc256[14:0]) ? cam_loc256 : 20'd0 ) |
 ( (snoop_in == cam_loc257[14:0]) ? cam_loc257 : 20'd0 ) |
 ( (snoop_in == cam_loc258[14:0]) ? cam_loc258 : 20'd0 ) |
 ( (snoop_in == cam_loc259[14:0]) ? cam_loc259 : 20'd0 ) |
 ( (snoop_in == cam_loc260[14:0]) ? cam_loc260 : 20'd0 ) |
 ( (snoop_in == cam_loc261[14:0]) ? cam_loc261 : 20'd0 ) |
 ( (snoop_in == cam_loc262[14:0]) ? cam_loc262 : 20'd0 ) |
 ( (snoop_in == cam_loc263[14:0]) ? cam_loc263 : 20'd0 ) |
 ( (snoop_in == cam_loc264[14:0]) ? cam_loc264 : 20'd0 ) |
 ( (snoop_in == cam_loc265[14:0]) ? cam_loc265 : 20'd0 ) |
 ( (snoop_in == cam_loc266[14:0]) ? cam_loc266 : 20'd0 ) |
 ( (snoop_in == cam_loc267[14:0]) ? cam_loc267 : 20'd0 ) |
 ( (snoop_in == cam_loc268[14:0]) ? cam_loc268 : 20'd0 ) |
 ( (snoop_in == cam_loc269[14:0]) ? cam_loc269 : 20'd0 ) |
 ( (snoop_in == cam_loc270[14:0]) ? cam_loc270 : 20'd0 ) |
 ( (snoop_in == cam_loc271[14:0]) ? cam_loc271 : 20'd0 ) |
 ( (snoop_in == cam_loc272[14:0]) ? cam_loc272 : 20'd0 ) |
 ( (snoop_in == cam_loc273[14:0]) ? cam_loc273 : 20'd0 ) |
 ( (snoop_in == cam_loc274[14:0]) ? cam_loc274 : 20'd0 ) |
 ( (snoop_in == cam_loc275[14:0]) ? cam_loc275 : 20'd0 ) |
 ( (snoop_in == cam_loc276[14:0]) ? cam_loc276 : 20'd0 ) |
 ( (snoop_in == cam_loc277[14:0]) ? cam_loc277 : 20'd0 ) |
 ( (snoop_in == cam_loc278[14:0]) ? cam_loc278 : 20'd0 ) |
 ( (snoop_in == cam_loc279[14:0]) ? cam_loc279 : 20'd0 ) |
 ( (snoop_in == cam_loc280[14:0]) ? cam_loc280 : 20'd0 ) |
 ( (snoop_in == cam_loc281[14:0]) ? cam_loc281 : 20'd0 ) |
 ( (snoop_in == cam_loc282[14:0]) ? cam_loc282 : 20'd0 ) |
 ( (snoop_in == cam_loc283[14:0]) ? cam_loc283 : 20'd0 ) |
 ( (snoop_in == cam_loc284[14:0]) ? cam_loc284 : 20'd0 ) |
 ( (snoop_in == cam_loc285[14:0]) ? cam_loc285 : 20'd0 ) |
 ( (snoop_in == cam_loc286[14:0]) ? cam_loc286 : 20'd0 ) |
 ( (snoop_in == cam_loc287[14:0]) ? cam_loc287 : 20'd0 ) |
 ( (snoop_in == cam_loc288[14:0]) ? cam_loc288 : 20'd0 ) |
 ( (snoop_in == cam_loc289[14:0]) ? cam_loc289 : 20'd0 ) |
 ( (snoop_in == cam_loc290[14:0]) ? cam_loc290 : 20'd0 ) |
 ( (snoop_in == cam_loc291[14:0]) ? cam_loc291 : 20'd0 ) |
 ( (snoop_in == cam_loc292[14:0]) ? cam_loc292 : 20'd0 ) |
 ( (snoop_in == cam_loc293[14:0]) ? cam_loc293 : 20'd0 ) |
 ( (snoop_in == cam_loc294[14:0]) ? cam_loc294 : 20'd0 ) |
 ( (snoop_in == cam_loc295[14:0]) ? cam_loc295 : 20'd0 ) |
 ( (snoop_in == cam_loc296[14:0]) ? cam_loc296 : 20'd0 ) |
 ( (snoop_in == cam_loc297[14:0]) ? cam_loc297 : 20'd0 ) |
 ( (snoop_in == cam_loc298[14:0]) ? cam_loc298 : 20'd0 ) |
 ( (snoop_in == cam_loc299[14:0]) ? cam_loc299 : 20'd0 ) |
 ( (snoop_in == cam_loc300[14:0]) ? cam_loc300 : 20'd0 ) |
 ( (snoop_in == cam_loc301[14:0]) ? cam_loc301 : 20'd0 ) |
 ( (snoop_in == cam_loc302[14:0]) ? cam_loc302 : 20'd0 ) |
 ( (snoop_in == cam_loc303[14:0]) ? cam_loc303 : 20'd0 ) |
 ( (snoop_in == cam_loc304[14:0]) ? cam_loc304 : 20'd0 ) |
 ( (snoop_in == cam_loc305[14:0]) ? cam_loc305 : 20'd0 ) |
 ( (snoop_in == cam_loc306[14:0]) ? cam_loc306 : 20'd0 ) |
 ( (snoop_in == cam_loc307[14:0]) ? cam_loc307 : 20'd0 ) |
 ( (snoop_in == cam_loc308[14:0]) ? cam_loc308 : 20'd0 ) |
 ( (snoop_in == cam_loc309[14:0]) ? cam_loc309 : 20'd0 ) |
 ( (snoop_in == cam_loc310[14:0]) ? cam_loc310 : 20'd0 ) |
 ( (snoop_in == cam_loc311[14:0]) ? cam_loc311 : 20'd0 ) |
 ( (snoop_in == cam_loc312[14:0]) ? cam_loc312 : 20'd0 ) |
 ( (snoop_in == cam_loc313[14:0]) ? cam_loc313 : 20'd0 ) |
 ( (snoop_in == cam_loc314[14:0]) ? cam_loc314 : 20'd0 ) |
 ( (snoop_in == cam_loc315[14:0]) ? cam_loc315 : 20'd0 ) |
 ( (snoop_in == cam_loc316[14:0]) ? cam_loc316 : 20'd0 ) |
 ( (snoop_in == cam_loc317[14:0]) ? cam_loc317 : 20'd0 ) |
 ( (snoop_in == cam_loc318[14:0]) ? cam_loc318 : 20'd0 ) |
 ( (snoop_in == cam_loc319[14:0]) ? cam_loc319 : 20'd0 ) |
 ( (snoop_in == cam_loc320[14:0]) ? cam_loc320 : 20'd0 ) |
 ( (snoop_in == cam_loc321[14:0]) ? cam_loc321 : 20'd0 ) |
 ( (snoop_in == cam_loc322[14:0]) ? cam_loc322 : 20'd0 ) |
 ( (snoop_in == cam_loc323[14:0]) ? cam_loc323 : 20'd0 ) |
 ( (snoop_in == cam_loc324[14:0]) ? cam_loc324 : 20'd0 ) |
 ( (snoop_in == cam_loc325[14:0]) ? cam_loc325 : 20'd0 ) |
 ( (snoop_in == cam_loc326[14:0]) ? cam_loc326 : 20'd0 ) |
 ( (snoop_in == cam_loc327[14:0]) ? cam_loc327 : 20'd0 ) |
 ( (snoop_in == cam_loc328[14:0]) ? cam_loc328 : 20'd0 ) |
 ( (snoop_in == cam_loc329[14:0]) ? cam_loc329 : 20'd0 ) |
 ( (snoop_in == cam_loc330[14:0]) ? cam_loc330 : 20'd0 ) |
 ( (snoop_in == cam_loc331[14:0]) ? cam_loc331 : 20'd0 ) |
 ( (snoop_in == cam_loc332[14:0]) ? cam_loc332 : 20'd0 ) |
 ( (snoop_in == cam_loc333[14:0]) ? cam_loc333 : 20'd0 ) |
 ( (snoop_in == cam_loc334[14:0]) ? cam_loc334 : 20'd0 ) |
 ( (snoop_in == cam_loc335[14:0]) ? cam_loc335 : 20'd0 ) |
 ( (snoop_in == cam_loc336[14:0]) ? cam_loc336 : 20'd0 ) |
 ( (snoop_in == cam_loc337[14:0]) ? cam_loc337 : 20'd0 ) |
 ( (snoop_in == cam_loc338[14:0]) ? cam_loc338 : 20'd0 ) |
 ( (snoop_in == cam_loc339[14:0]) ? cam_loc339 : 20'd0 ) |
 ( (snoop_in == cam_loc340[14:0]) ? cam_loc340 : 20'd0 ) |
 ( (snoop_in == cam_loc341[14:0]) ? cam_loc341 : 20'd0 ) |
 ( (snoop_in == cam_loc342[14:0]) ? cam_loc342 : 20'd0 ) |
 ( (snoop_in == cam_loc343[14:0]) ? cam_loc343 : 20'd0 ) |
 ( (snoop_in == cam_loc344[14:0]) ? cam_loc344 : 20'd0 ) |
 ( (snoop_in == cam_loc345[14:0]) ? cam_loc345 : 20'd0 ) |
 ( (snoop_in == cam_loc346[14:0]) ? cam_loc346 : 20'd0 ) |
 ( (snoop_in == cam_loc347[14:0]) ? cam_loc347 : 20'd0 ) |
 ( (snoop_in == cam_loc348[14:0]) ? cam_loc348 : 20'd0 ) |
 ( (snoop_in == cam_loc349[14:0]) ? cam_loc349 : 20'd0 ) |
 ( (snoop_in == cam_loc350[14:0]) ? cam_loc350 : 20'd0 ) |
 ( (snoop_in == cam_loc351[14:0]) ? cam_loc351 : 20'd0 ) |
 ( (snoop_in == cam_loc352[14:0]) ? cam_loc352 : 20'd0 ) |
 ( (snoop_in == cam_loc353[14:0]) ? cam_loc353 : 20'd0 ) |
 ( (snoop_in == cam_loc354[14:0]) ? cam_loc354 : 20'd0 ) |
 ( (snoop_in == cam_loc355[14:0]) ? cam_loc355 : 20'd0 ) |
 ( (snoop_in == cam_loc356[14:0]) ? cam_loc356 : 20'd0 ) |
 ( (snoop_in == cam_loc357[14:0]) ? cam_loc357 : 20'd0 ) |
 ( (snoop_in == cam_loc358[14:0]) ? cam_loc358 : 20'd0 ) |
 ( (snoop_in == cam_loc359[14:0]) ? cam_loc359 : 20'd0 ) |
 ( (snoop_in == cam_loc360[14:0]) ? cam_loc360 : 20'd0 ) |
 ( (snoop_in == cam_loc361[14:0]) ? cam_loc361 : 20'd0 ) |
 ( (snoop_in == cam_loc362[14:0]) ? cam_loc362 : 20'd0 ) |
 ( (snoop_in == cam_loc363[14:0]) ? cam_loc363 : 20'd0 ) |
 ( (snoop_in == cam_loc364[14:0]) ? cam_loc364 : 20'd0 ) |
 ( (snoop_in == cam_loc365[14:0]) ? cam_loc365 : 20'd0 ) |
 ( (snoop_in == cam_loc366[14:0]) ? cam_loc366 : 20'd0 ) |
 ( (snoop_in == cam_loc367[14:0]) ? cam_loc367 : 20'd0 ) |
 ( (snoop_in == cam_loc368[14:0]) ? cam_loc368 : 20'd0 ) |
 ( (snoop_in == cam_loc369[14:0]) ? cam_loc369 : 20'd0 ) |
 ( (snoop_in == cam_loc370[14:0]) ? cam_loc370 : 20'd0 ) |
 ( (snoop_in == cam_loc371[14:0]) ? cam_loc371 : 20'd0 ) |
 ( (snoop_in == cam_loc372[14:0]) ? cam_loc372 : 20'd0 ) |
 ( (snoop_in == cam_loc373[14:0]) ? cam_loc373 : 20'd0 ) |
 ( (snoop_in == cam_loc374[14:0]) ? cam_loc374 : 20'd0 ) |
 ( (snoop_in == cam_loc375[14:0]) ? cam_loc375 : 20'd0 ) |
 ( (snoop_in == cam_loc376[14:0]) ? cam_loc376 : 20'd0 ) |
 ( (snoop_in == cam_loc377[14:0]) ? cam_loc377 : 20'd0 ) |
 ( (snoop_in == cam_loc378[14:0]) ? cam_loc378 : 20'd0 ) |
 ( (snoop_in == cam_loc379[14:0]) ? cam_loc379 : 20'd0 ) |
 ( (snoop_in == cam_loc380[14:0]) ? cam_loc380 : 20'd0 ) |
 ( (snoop_in == cam_loc381[14:0]) ? cam_loc381 : 20'd0 ) |
 ( (snoop_in == cam_loc382[14:0]) ? cam_loc382 : 20'd0 ) |
 ( (snoop_in == cam_loc383[14:0]) ? cam_loc383 : 20'd0 ) |
 ( (snoop_in == cam_loc384[14:0]) ? cam_loc384 : 20'd0 ) |
 ( (snoop_in == cam_loc385[14:0]) ? cam_loc385 : 20'd0 ) |
 ( (snoop_in == cam_loc386[14:0]) ? cam_loc386 : 20'd0 ) |
 ( (snoop_in == cam_loc387[14:0]) ? cam_loc387 : 20'd0 ) |
 ( (snoop_in == cam_loc388[14:0]) ? cam_loc388 : 20'd0 ) |
 ( (snoop_in == cam_loc389[14:0]) ? cam_loc389 : 20'd0 ) |
 ( (snoop_in == cam_loc390[14:0]) ? cam_loc390 : 20'd0 ) |
 ( (snoop_in == cam_loc391[14:0]) ? cam_loc391 : 20'd0 ) |
 ( (snoop_in == cam_loc392[14:0]) ? cam_loc392 : 20'd0 ) |
 ( (snoop_in == cam_loc393[14:0]) ? cam_loc393 : 20'd0 ) |
 ( (snoop_in == cam_loc394[14:0]) ? cam_loc394 : 20'd0 ) |
 ( (snoop_in == cam_loc395[14:0]) ? cam_loc395 : 20'd0 ) |
 ( (snoop_in == cam_loc396[14:0]) ? cam_loc396 : 20'd0 ) |
 ( (snoop_in == cam_loc397[14:0]) ? cam_loc397 : 20'd0 ) |
 ( (snoop_in == cam_loc398[14:0]) ? cam_loc398 : 20'd0 ) |
 ( (snoop_in == cam_loc399[14:0]) ? cam_loc399 : 20'd0 ) |
 ( (snoop_in == cam_loc400[14:0]) ? cam_loc400 : 20'd0 ) |
 ( (snoop_in == cam_loc401[14:0]) ? cam_loc401 : 20'd0 ) |
 ( (snoop_in == cam_loc402[14:0]) ? cam_loc402 : 20'd0 ) |
 ( (snoop_in == cam_loc403[14:0]) ? cam_loc403 : 20'd0 ) |
 ( (snoop_in == cam_loc404[14:0]) ? cam_loc404 : 20'd0 ) |
 ( (snoop_in == cam_loc405[14:0]) ? cam_loc405 : 20'd0 ) |
 ( (snoop_in == cam_loc406[14:0]) ? cam_loc406 : 20'd0 ) |
 ( (snoop_in == cam_loc407[14:0]) ? cam_loc407 : 20'd0 ) |
 ( (snoop_in == cam_loc408[14:0]) ? cam_loc408 : 20'd0 ) |
 ( (snoop_in == cam_loc409[14:0]) ? cam_loc409 : 20'd0 ) |
 ( (snoop_in == cam_loc410[14:0]) ? cam_loc410 : 20'd0 ) |
 ( (snoop_in == cam_loc411[14:0]) ? cam_loc411 : 20'd0 ) |
 ( (snoop_in == cam_loc412[14:0]) ? cam_loc412 : 20'd0 ) |
 ( (snoop_in == cam_loc413[14:0]) ? cam_loc413 : 20'd0 ) |
 ( (snoop_in == cam_loc414[14:0]) ? cam_loc414 : 20'd0 ) |
 ( (snoop_in == cam_loc415[14:0]) ? cam_loc415 : 20'd0 ) |
 ( (snoop_in == cam_loc416[14:0]) ? cam_loc416 : 20'd0 ) |
 ( (snoop_in == cam_loc417[14:0]) ? cam_loc417 : 20'd0 ) |
 ( (snoop_in == cam_loc418[14:0]) ? cam_loc418 : 20'd0 ) |
 ( (snoop_in == cam_loc419[14:0]) ? cam_loc419 : 20'd0 ) |
 ( (snoop_in == cam_loc420[14:0]) ? cam_loc420 : 20'd0 ) |
 ( (snoop_in == cam_loc421[14:0]) ? cam_loc421 : 20'd0 ) |
 ( (snoop_in == cam_loc422[14:0]) ? cam_loc422 : 20'd0 ) |
 ( (snoop_in == cam_loc423[14:0]) ? cam_loc423 : 20'd0 ) |
 ( (snoop_in == cam_loc424[14:0]) ? cam_loc424 : 20'd0 ) |
 ( (snoop_in == cam_loc425[14:0]) ? cam_loc425 : 20'd0 ) |
 ( (snoop_in == cam_loc426[14:0]) ? cam_loc426 : 20'd0 ) |
 ( (snoop_in == cam_loc427[14:0]) ? cam_loc427 : 20'd0 ) |
 ( (snoop_in == cam_loc428[14:0]) ? cam_loc428 : 20'd0 ) |
 ( (snoop_in == cam_loc429[14:0]) ? cam_loc429 : 20'd0 ) |
 ( (snoop_in == cam_loc430[14:0]) ? cam_loc430 : 20'd0 ) |
 ( (snoop_in == cam_loc431[14:0]) ? cam_loc431 : 20'd0 ) |
 ( (snoop_in == cam_loc432[14:0]) ? cam_loc432 : 20'd0 ) |
 ( (snoop_in == cam_loc433[14:0]) ? cam_loc433 : 20'd0 ) |
 ( (snoop_in == cam_loc434[14:0]) ? cam_loc434 : 20'd0 ) |
 ( (snoop_in == cam_loc435[14:0]) ? cam_loc435 : 20'd0 ) |
 ( (snoop_in == cam_loc436[14:0]) ? cam_loc436 : 20'd0 ) |
 ( (snoop_in == cam_loc437[14:0]) ? cam_loc437 : 20'd0 ) |
 ( (snoop_in == cam_loc438[14:0]) ? cam_loc438 : 20'd0 ) |
 ( (snoop_in == cam_loc439[14:0]) ? cam_loc439 : 20'd0 ) |
 ( (snoop_in == cam_loc440[14:0]) ? cam_loc440 : 20'd0 ) |
 ( (snoop_in == cam_loc441[14:0]) ? cam_loc441 : 20'd0 ) |
 ( (snoop_in == cam_loc442[14:0]) ? cam_loc442 : 20'd0 ) |
 ( (snoop_in == cam_loc443[14:0]) ? cam_loc443 : 20'd0 ) |
 ( (snoop_in == cam_loc444[14:0]) ? cam_loc444 : 20'd0 ) |
 ( (snoop_in == cam_loc445[14:0]) ? cam_loc445 : 20'd0 ) |
 ( (snoop_in == cam_loc446[14:0]) ? cam_loc446 : 20'd0 ) |
 ( (snoop_in == cam_loc447[14:0]) ? cam_loc447 : 20'd0 ) |
 ( (snoop_in == cam_loc448[14:0]) ? cam_loc448 : 20'd0 ) |
 ( (snoop_in == cam_loc449[14:0]) ? cam_loc449 : 20'd0 ) |
 ( (snoop_in == cam_loc450[14:0]) ? cam_loc450 : 20'd0 ) |
 ( (snoop_in == cam_loc451[14:0]) ? cam_loc451 : 20'd0 ) |
 ( (snoop_in == cam_loc452[14:0]) ? cam_loc452 : 20'd0 ) |
 ( (snoop_in == cam_loc453[14:0]) ? cam_loc453 : 20'd0 ) |
 ( (snoop_in == cam_loc454[14:0]) ? cam_loc454 : 20'd0 ) |
 ( (snoop_in == cam_loc455[14:0]) ? cam_loc455 : 20'd0 ) |
 ( (snoop_in == cam_loc456[14:0]) ? cam_loc456 : 20'd0 ) |
 ( (snoop_in == cam_loc457[14:0]) ? cam_loc457 : 20'd0 ) |
 ( (snoop_in == cam_loc458[14:0]) ? cam_loc458 : 20'd0 ) |
 ( (snoop_in == cam_loc459[14:0]) ? cam_loc459 : 20'd0 ) |
 ( (snoop_in == cam_loc460[14:0]) ? cam_loc460 : 20'd0 ) |
 ( (snoop_in == cam_loc461[14:0]) ? cam_loc461 : 20'd0 ) |
 ( (snoop_in == cam_loc462[14:0]) ? cam_loc462 : 20'd0 ) |
 ( (snoop_in == cam_loc463[14:0]) ? cam_loc463 : 20'd0 ) |
 ( (snoop_in == cam_loc464[14:0]) ? cam_loc464 : 20'd0 ) |
 ( (snoop_in == cam_loc465[14:0]) ? cam_loc465 : 20'd0 ) |
 ( (snoop_in == cam_loc466[14:0]) ? cam_loc466 : 20'd0 ) |
 ( (snoop_in == cam_loc467[14:0]) ? cam_loc467 : 20'd0 ) |
 ( (snoop_in == cam_loc468[14:0]) ? cam_loc468 : 20'd0 ) |
 ( (snoop_in == cam_loc469[14:0]) ? cam_loc469 : 20'd0 ) |
 ( (snoop_in == cam_loc470[14:0]) ? cam_loc470 : 20'd0 ) |
 ( (snoop_in == cam_loc471[14:0]) ? cam_loc471 : 20'd0 ) |
 ( (snoop_in == cam_loc472[14:0]) ? cam_loc472 : 20'd0 ) |
 ( (snoop_in == cam_loc473[14:0]) ? cam_loc473 : 20'd0 ) |
 ( (snoop_in == cam_loc474[14:0]) ? cam_loc474 : 20'd0 ) |
 ( (snoop_in == cam_loc475[14:0]) ? cam_loc475 : 20'd0 ) |
 ( (snoop_in == cam_loc476[14:0]) ? cam_loc476 : 20'd0 ) |
 ( (snoop_in == cam_loc477[14:0]) ? cam_loc477 : 20'd0 ) |
 ( (snoop_in == cam_loc478[14:0]) ? cam_loc478 : 20'd0 ) |
 ( (snoop_in == cam_loc479[14:0]) ? cam_loc479 : 20'd0 ) |
 ( (snoop_in == cam_loc480[14:0]) ? cam_loc480 : 20'd0 ) |
 ( (snoop_in == cam_loc481[14:0]) ? cam_loc481 : 20'd0 ) |
 ( (snoop_in == cam_loc482[14:0]) ? cam_loc482 : 20'd0 ) |
 ( (snoop_in == cam_loc483[14:0]) ? cam_loc483 : 20'd0 ) |
 ( (snoop_in == cam_loc484[14:0]) ? cam_loc484 : 20'd0 ) |
 ( (snoop_in == cam_loc485[14:0]) ? cam_loc485 : 20'd0 ) |
 ( (snoop_in == cam_loc486[14:0]) ? cam_loc486 : 20'd0 ) |
 ( (snoop_in == cam_loc487[14:0]) ? cam_loc487 : 20'd0 ) |
 ( (snoop_in == cam_loc488[14:0]) ? cam_loc488 : 20'd0 ) |
 ( (snoop_in == cam_loc489[14:0]) ? cam_loc489 : 20'd0 ) |
 ( (snoop_in == cam_loc490[14:0]) ? cam_loc490 : 20'd0 ) |
 ( (snoop_in == cam_loc491[14:0]) ? cam_loc491 : 20'd0 ) |
 ( (snoop_in == cam_loc492[14:0]) ? cam_loc492 : 20'd0 ) |
 ( (snoop_in == cam_loc493[14:0]) ? cam_loc493 : 20'd0 ) |
 ( (snoop_in == cam_loc494[14:0]) ? cam_loc494 : 20'd0 ) |
 ( (snoop_in == cam_loc495[14:0]) ? cam_loc495 : 20'd0 ) |
 ( (snoop_in == cam_loc496[14:0]) ? cam_loc496 : 20'd0 ) |
 ( (snoop_in == cam_loc497[14:0]) ? cam_loc497 : 20'd0 ) |
 ( (snoop_in == cam_loc498[14:0]) ? cam_loc498 : 20'd0 ) |
 ( (snoop_in == cam_loc499[14:0]) ? cam_loc499 : 20'd0 ) |
 ( (snoop_in == cam_loc500[14:0]) ? cam_loc500 : 20'd0 ) |
 ( (snoop_in == cam_loc501[14:0]) ? cam_loc501 : 20'd0 ) |
 ( (snoop_in == cam_loc502[14:0]) ? cam_loc502 : 20'd0 ) |
 ( (snoop_in == cam_loc503[14:0]) ? cam_loc503 : 20'd0 ) |
 ( (snoop_in == cam_loc504[14:0]) ? cam_loc504 : 20'd0 ) |
 ( (snoop_in == cam_loc505[14:0]) ? cam_loc505 : 20'd0 ) |
 ( (snoop_in == cam_loc506[14:0]) ? cam_loc506 : 20'd0 ) |
 ( (snoop_in == cam_loc507[14:0]) ? cam_loc507 : 20'd0 ) |
 ( (snoop_in == cam_loc508[14:0]) ? cam_loc508 : 20'd0 ) |
 ( (snoop_in == cam_loc509[14:0]) ? cam_loc509 : 20'd0 ) |
 ( (snoop_in == cam_loc510[14:0]) ? cam_loc510 : 20'd0 ) |
 ( (snoop_in == cam_loc511[14:0]) ? cam_loc511 : 20'd0 ) |
 ( (snoop_in == cam_loc512[14:0]) ? cam_loc512 : 20'd0 ) |
 ( (snoop_in == cam_loc513[14:0]) ? cam_loc513 : 20'd0 ) |
 ( (snoop_in == cam_loc514[14:0]) ? cam_loc514 : 20'd0 ) |
 ( (snoop_in == cam_loc515[14:0]) ? cam_loc515 : 20'd0 ) |
 ( (snoop_in == cam_loc516[14:0]) ? cam_loc516 : 20'd0 ) |
 ( (snoop_in == cam_loc517[14:0]) ? cam_loc517 : 20'd0 ) |
 ( (snoop_in == cam_loc518[14:0]) ? cam_loc518 : 20'd0 ) |
 ( (snoop_in == cam_loc519[14:0]) ? cam_loc519 : 20'd0 ) |
 ( (snoop_in == cam_loc520[14:0]) ? cam_loc520 : 20'd0 ) |
 ( (snoop_in == cam_loc521[14:0]) ? cam_loc521 : 20'd0 ) |
 ( (snoop_in == cam_loc522[14:0]) ? cam_loc522 : 20'd0 ) |
 ( (snoop_in == cam_loc523[14:0]) ? cam_loc523 : 20'd0 ) |
 ( (snoop_in == cam_loc524[14:0]) ? cam_loc524 : 20'd0 ) |
 ( (snoop_in == cam_loc525[14:0]) ? cam_loc525 : 20'd0 ) |
 ( (snoop_in == cam_loc526[14:0]) ? cam_loc526 : 20'd0 ) |
 ( (snoop_in == cam_loc527[14:0]) ? cam_loc527 : 20'd0 ) |
 ( (snoop_in == cam_loc528[14:0]) ? cam_loc528 : 20'd0 ) |
 ( (snoop_in == cam_loc529[14:0]) ? cam_loc529 : 20'd0 ) |
 ( (snoop_in == cam_loc530[14:0]) ? cam_loc530 : 20'd0 ) |
 ( (snoop_in == cam_loc531[14:0]) ? cam_loc531 : 20'd0 ) |
 ( (snoop_in == cam_loc532[14:0]) ? cam_loc532 : 20'd0 ) |
 ( (snoop_in == cam_loc533[14:0]) ? cam_loc533 : 20'd0 ) |
 ( (snoop_in == cam_loc534[14:0]) ? cam_loc534 : 20'd0 ) |
 ( (snoop_in == cam_loc535[14:0]) ? cam_loc535 : 20'd0 ) |
 ( (snoop_in == cam_loc536[14:0]) ? cam_loc536 : 20'd0 ) |
 ( (snoop_in == cam_loc537[14:0]) ? cam_loc537 : 20'd0 ) |
 ( (snoop_in == cam_loc538[14:0]) ? cam_loc538 : 20'd0 ) |
 ( (snoop_in == cam_loc539[14:0]) ? cam_loc539 : 20'd0 ) |
 ( (snoop_in == cam_loc540[14:0]) ? cam_loc540 : 20'd0 ) |
 ( (snoop_in == cam_loc541[14:0]) ? cam_loc541 : 20'd0 ) |
 ( (snoop_in == cam_loc542[14:0]) ? cam_loc542 : 20'd0 ) |
 ( (snoop_in == cam_loc543[14:0]) ? cam_loc543 : 20'd0 ) |
 ( (snoop_in == cam_loc544[14:0]) ? cam_loc544 : 20'd0 ) |
 ( (snoop_in == cam_loc545[14:0]) ? cam_loc545 : 20'd0 ) |
 ( (snoop_in == cam_loc546[14:0]) ? cam_loc546 : 20'd0 ) |
 ( (snoop_in == cam_loc547[14:0]) ? cam_loc547 : 20'd0 ) |
 ( (snoop_in == cam_loc548[14:0]) ? cam_loc548 : 20'd0 ) |
 ( (snoop_in == cam_loc549[14:0]) ? cam_loc549 : 20'd0 ) |
 ( (snoop_in == cam_loc550[14:0]) ? cam_loc550 : 20'd0 ) |
 ( (snoop_in == cam_loc551[14:0]) ? cam_loc551 : 20'd0 ) |
 ( (snoop_in == cam_loc552[14:0]) ? cam_loc552 : 20'd0 ) |
 ( (snoop_in == cam_loc553[14:0]) ? cam_loc553 : 20'd0 ) |
 ( (snoop_in == cam_loc554[14:0]) ? cam_loc554 : 20'd0 ) |
 ( (snoop_in == cam_loc555[14:0]) ? cam_loc555 : 20'd0 ) |
 ( (snoop_in == cam_loc556[14:0]) ? cam_loc556 : 20'd0 ) |
 ( (snoop_in == cam_loc557[14:0]) ? cam_loc557 : 20'd0 ) |
 ( (snoop_in == cam_loc558[14:0]) ? cam_loc558 : 20'd0 ) |
 ( (snoop_in == cam_loc559[14:0]) ? cam_loc559 : 20'd0 ) |
 ( (snoop_in == cam_loc560[14:0]) ? cam_loc560 : 20'd0 ) |
 ( (snoop_in == cam_loc561[14:0]) ? cam_loc561 : 20'd0 ) |
 ( (snoop_in == cam_loc562[14:0]) ? cam_loc562 : 20'd0 ) |
 ( (snoop_in == cam_loc563[14:0]) ? cam_loc563 : 20'd0 ) |
 ( (snoop_in == cam_loc564[14:0]) ? cam_loc564 : 20'd0 ) |
 ( (snoop_in == cam_loc565[14:0]) ? cam_loc565 : 20'd0 ) |
 ( (snoop_in == cam_loc566[14:0]) ? cam_loc566 : 20'd0 ) |
 ( (snoop_in == cam_loc567[14:0]) ? cam_loc567 : 20'd0 ) |
 ( (snoop_in == cam_loc568[14:0]) ? cam_loc568 : 20'd0 ) |
 ( (snoop_in == cam_loc569[14:0]) ? cam_loc569 : 20'd0 ) |
 ( (snoop_in == cam_loc570[14:0]) ? cam_loc570 : 20'd0 ) |
 ( (snoop_in == cam_loc571[14:0]) ? cam_loc571 : 20'd0 ) |
 ( (snoop_in == cam_loc572[14:0]) ? cam_loc572 : 20'd0 ) |
 ( (snoop_in == cam_loc573[14:0]) ? cam_loc573 : 20'd0 ) |
 ( (snoop_in == cam_loc574[14:0]) ? cam_loc574 : 20'd0 ) |
 ( (snoop_in == cam_loc575[14:0]) ? cam_loc575 : 20'd0 ) |
 ( (snoop_in == cam_loc576[14:0]) ? cam_loc576 : 20'd0 ) |
 ( (snoop_in == cam_loc577[14:0]) ? cam_loc577 : 20'd0 ) |
 ( (snoop_in == cam_loc578[14:0]) ? cam_loc578 : 20'd0 ) |
 ( (snoop_in == cam_loc579[14:0]) ? cam_loc579 : 20'd0 ) |
 ( (snoop_in == cam_loc580[14:0]) ? cam_loc580 : 20'd0 ) |
 ( (snoop_in == cam_loc581[14:0]) ? cam_loc581 : 20'd0 ) |
 ( (snoop_in == cam_loc582[14:0]) ? cam_loc582 : 20'd0 ) |
 ( (snoop_in == cam_loc583[14:0]) ? cam_loc583 : 20'd0 ) |
 ( (snoop_in == cam_loc584[14:0]) ? cam_loc584 : 20'd0 ) |
 ( (snoop_in == cam_loc585[14:0]) ? cam_loc585 : 20'd0 ) |
 ( (snoop_in == cam_loc586[14:0]) ? cam_loc586 : 20'd0 ) |
 ( (snoop_in == cam_loc587[14:0]) ? cam_loc587 : 20'd0 ) |
 ( (snoop_in == cam_loc588[14:0]) ? cam_loc588 : 20'd0 ) |
 ( (snoop_in == cam_loc589[14:0]) ? cam_loc589 : 20'd0 ) |
 ( (snoop_in == cam_loc590[14:0]) ? cam_loc590 : 20'd0 ) |
 ( (snoop_in == cam_loc591[14:0]) ? cam_loc591 : 20'd0 ) |
 ( (snoop_in == cam_loc592[14:0]) ? cam_loc592 : 20'd0 ) |
 ( (snoop_in == cam_loc593[14:0]) ? cam_loc593 : 20'd0 ) |
 ( (snoop_in == cam_loc594[14:0]) ? cam_loc594 : 20'd0 ) |
 ( (snoop_in == cam_loc595[14:0]) ? cam_loc595 : 20'd0 ) |
 ( (snoop_in == cam_loc596[14:0]) ? cam_loc596 : 20'd0 ) |
 ( (snoop_in == cam_loc597[14:0]) ? cam_loc597 : 20'd0 ) |
 ( (snoop_in == cam_loc598[14:0]) ? cam_loc598 : 20'd0 ) |
 ( (snoop_in == cam_loc599[14:0]) ? cam_loc599 : 20'd0 ) |
 ( (snoop_in == cam_loc600[14:0]) ? cam_loc600 : 20'd0 ) |
 ( (snoop_in == cam_loc601[14:0]) ? cam_loc601 : 20'd0 ) |
 ( (snoop_in == cam_loc602[14:0]) ? cam_loc602 : 20'd0 ) |
 ( (snoop_in == cam_loc603[14:0]) ? cam_loc603 : 20'd0 ) |
 ( (snoop_in == cam_loc604[14:0]) ? cam_loc604 : 20'd0 ) |
 ( (snoop_in == cam_loc605[14:0]) ? cam_loc605 : 20'd0 ) |
 ( (snoop_in == cam_loc606[14:0]) ? cam_loc606 : 20'd0 ) |
 ( (snoop_in == cam_loc607[14:0]) ? cam_loc607 : 20'd0 ) |
 ( (snoop_in == cam_loc608[14:0]) ? cam_loc608 : 20'd0 ) |
 ( (snoop_in == cam_loc609[14:0]) ? cam_loc609 : 20'd0 ) |
 ( (snoop_in == cam_loc610[14:0]) ? cam_loc610 : 20'd0 ) |
 ( (snoop_in == cam_loc611[14:0]) ? cam_loc611 : 20'd0 ) |
 ( (snoop_in == cam_loc612[14:0]) ? cam_loc612 : 20'd0 ) |
 ( (snoop_in == cam_loc613[14:0]) ? cam_loc613 : 20'd0 ) |
 ( (snoop_in == cam_loc614[14:0]) ? cam_loc614 : 20'd0 ) |
 ( (snoop_in == cam_loc615[14:0]) ? cam_loc615 : 20'd0 ) |
 ( (snoop_in == cam_loc616[14:0]) ? cam_loc616 : 20'd0 ) |
 ( (snoop_in == cam_loc617[14:0]) ? cam_loc617 : 20'd0 ) |
 ( (snoop_in == cam_loc618[14:0]) ? cam_loc618 : 20'd0 ) |
 ( (snoop_in == cam_loc619[14:0]) ? cam_loc619 : 20'd0 ) |
 ( (snoop_in == cam_loc620[14:0]) ? cam_loc620 : 20'd0 ) |
 ( (snoop_in == cam_loc621[14:0]) ? cam_loc621 : 20'd0 ) |
 ( (snoop_in == cam_loc622[14:0]) ? cam_loc622 : 20'd0 ) |
 ( (snoop_in == cam_loc623[14:0]) ? cam_loc623 : 20'd0 ) |
 ( (snoop_in == cam_loc624[14:0]) ? cam_loc624 : 20'd0 ) |
 ( (snoop_in == cam_loc625[14:0]) ? cam_loc625 : 20'd0 ) |
 ( (snoop_in == cam_loc626[14:0]) ? cam_loc626 : 20'd0 ) |
 ( (snoop_in == cam_loc627[14:0]) ? cam_loc627 : 20'd0 ) |
 ( (snoop_in == cam_loc628[14:0]) ? cam_loc628 : 20'd0 ) |
 ( (snoop_in == cam_loc629[14:0]) ? cam_loc629 : 20'd0 ) |
 ( (snoop_in == cam_loc630[14:0]) ? cam_loc630 : 20'd0 ) |
 ( (snoop_in == cam_loc631[14:0]) ? cam_loc631 : 20'd0 ) |
 ( (snoop_in == cam_loc632[14:0]) ? cam_loc632 : 20'd0 ) |
 ( (snoop_in == cam_loc633[14:0]) ? cam_loc633 : 20'd0 ) |
 ( (snoop_in == cam_loc634[14:0]) ? cam_loc634 : 20'd0 ) |
 ( (snoop_in == cam_loc635[14:0]) ? cam_loc635 : 20'd0 ) |
 ( (snoop_in == cam_loc636[14:0]) ? cam_loc636 : 20'd0 ) |
 ( (snoop_in == cam_loc637[14:0]) ? cam_loc637 : 20'd0 ) |
 ( (snoop_in == cam_loc638[14:0]) ? cam_loc638 : 20'd0 ) |
 ( (snoop_in == cam_loc639[14:0]) ? cam_loc639 : 20'd0 ) |
 ( (snoop_in == cam_loc640[14:0]) ? cam_loc640 : 20'd0 ) |
 ( (snoop_in == cam_loc641[14:0]) ? cam_loc641 : 20'd0 ) |
 ( (snoop_in == cam_loc642[14:0]) ? cam_loc642 : 20'd0 ) |
 ( (snoop_in == cam_loc643[14:0]) ? cam_loc643 : 20'd0 ) |
 ( (snoop_in == cam_loc644[14:0]) ? cam_loc644 : 20'd0 ) |
 ( (snoop_in == cam_loc645[14:0]) ? cam_loc645 : 20'd0 ) |
 ( (snoop_in == cam_loc646[14:0]) ? cam_loc646 : 20'd0 ) |
 ( (snoop_in == cam_loc647[14:0]) ? cam_loc647 : 20'd0 ) |
 ( (snoop_in == cam_loc648[14:0]) ? cam_loc648 : 20'd0 ) |
 ( (snoop_in == cam_loc649[14:0]) ? cam_loc649 : 20'd0 ) |
 ( (snoop_in == cam_loc650[14:0]) ? cam_loc650 : 20'd0 ) |
 ( (snoop_in == cam_loc651[14:0]) ? cam_loc651 : 20'd0 ) |
 ( (snoop_in == cam_loc652[14:0]) ? cam_loc652 : 20'd0 ) |
 ( (snoop_in == cam_loc653[14:0]) ? cam_loc653 : 20'd0 ) |
 ( (snoop_in == cam_loc654[14:0]) ? cam_loc654 : 20'd0 ) |
 ( (snoop_in == cam_loc655[14:0]) ? cam_loc655 : 20'd0 ) |
 ( (snoop_in == cam_loc656[14:0]) ? cam_loc656 : 20'd0 ) |
 ( (snoop_in == cam_loc657[14:0]) ? cam_loc657 : 20'd0 ) |
 ( (snoop_in == cam_loc658[14:0]) ? cam_loc658 : 20'd0 ) |
 ( (snoop_in == cam_loc659[14:0]) ? cam_loc659 : 20'd0 ) |
 ( (snoop_in == cam_loc660[14:0]) ? cam_loc660 : 20'd0 ) |
 ( (snoop_in == cam_loc661[14:0]) ? cam_loc661 : 20'd0 ) |
 ( (snoop_in == cam_loc662[14:0]) ? cam_loc662 : 20'd0 ) |
 ( (snoop_in == cam_loc663[14:0]) ? cam_loc663 : 20'd0 ) |
 ( (snoop_in == cam_loc664[14:0]) ? cam_loc664 : 20'd0 ) |
 ( (snoop_in == cam_loc665[14:0]) ? cam_loc665 : 20'd0 ) |
 ( (snoop_in == cam_loc666[14:0]) ? cam_loc666 : 20'd0 ) |
 ( (snoop_in == cam_loc667[14:0]) ? cam_loc667 : 20'd0 ) |
 ( (snoop_in == cam_loc668[14:0]) ? cam_loc668 : 20'd0 ) |
 ( (snoop_in == cam_loc669[14:0]) ? cam_loc669 : 20'd0 ) |
 ( (snoop_in == cam_loc670[14:0]) ? cam_loc670 : 20'd0 ) |
 ( (snoop_in == cam_loc671[14:0]) ? cam_loc671 : 20'd0 ) |
 ( (snoop_in == cam_loc672[14:0]) ? cam_loc672 : 20'd0 ) |
 ( (snoop_in == cam_loc673[14:0]) ? cam_loc673 : 20'd0 ) |
 ( (snoop_in == cam_loc674[14:0]) ? cam_loc674 : 20'd0 ) |
 ( (snoop_in == cam_loc675[14:0]) ? cam_loc675 : 20'd0 ) |
 ( (snoop_in == cam_loc676[14:0]) ? cam_loc676 : 20'd0 ) |
 ( (snoop_in == cam_loc677[14:0]) ? cam_loc677 : 20'd0 ) |
 ( (snoop_in == cam_loc678[14:0]) ? cam_loc678 : 20'd0 ) |
 ( (snoop_in == cam_loc679[14:0]) ? cam_loc679 : 20'd0 ) |
 ( (snoop_in == cam_loc680[14:0]) ? cam_loc680 : 20'd0 ) |
 ( (snoop_in == cam_loc681[14:0]) ? cam_loc681 : 20'd0 ) |
 ( (snoop_in == cam_loc682[14:0]) ? cam_loc682 : 20'd0 ) |
 ( (snoop_in == cam_loc683[14:0]) ? cam_loc683 : 20'd0 ) |
 ( (snoop_in == cam_loc684[14:0]) ? cam_loc684 : 20'd0 ) |
 ( (snoop_in == cam_loc685[14:0]) ? cam_loc685 : 20'd0 ) |
 ( (snoop_in == cam_loc686[14:0]) ? cam_loc686 : 20'd0 ) |
 ( (snoop_in == cam_loc687[14:0]) ? cam_loc687 : 20'd0 ) |
 ( (snoop_in == cam_loc688[14:0]) ? cam_loc688 : 20'd0 ) |
 ( (snoop_in == cam_loc689[14:0]) ? cam_loc689 : 20'd0 ) |
 ( (snoop_in == cam_loc690[14:0]) ? cam_loc690 : 20'd0 ) |
 ( (snoop_in == cam_loc691[14:0]) ? cam_loc691 : 20'd0 ) |
 ( (snoop_in == cam_loc692[14:0]) ? cam_loc692 : 20'd0 ) |
 ( (snoop_in == cam_loc693[14:0]) ? cam_loc693 : 20'd0 ) |
 ( (snoop_in == cam_loc694[14:0]) ? cam_loc694 : 20'd0 ) |
 ( (snoop_in == cam_loc695[14:0]) ? cam_loc695 : 20'd0 ) |
 ( (snoop_in == cam_loc696[14:0]) ? cam_loc696 : 20'd0 ) |
 ( (snoop_in == cam_loc697[14:0]) ? cam_loc697 : 20'd0 ) |
 ( (snoop_in == cam_loc698[14:0]) ? cam_loc698 : 20'd0 ) |
 ( (snoop_in == cam_loc699[14:0]) ? cam_loc699 : 20'd0 ) |
 ( (snoop_in == cam_loc700[14:0]) ? cam_loc700 : 20'd0 ) |
 ( (snoop_in == cam_loc701[14:0]) ? cam_loc701 : 20'd0 ) |
 ( (snoop_in == cam_loc702[14:0]) ? cam_loc702 : 20'd0 ) |
 ( (snoop_in == cam_loc703[14:0]) ? cam_loc703 : 20'd0 ) |
 ( (snoop_in == cam_loc704[14:0]) ? cam_loc704 : 20'd0 ) |
 ( (snoop_in == cam_loc705[14:0]) ? cam_loc705 : 20'd0 ) |
 ( (snoop_in == cam_loc706[14:0]) ? cam_loc706 : 20'd0 ) |
 ( (snoop_in == cam_loc707[14:0]) ? cam_loc707 : 20'd0 ) |
 ( (snoop_in == cam_loc708[14:0]) ? cam_loc708 : 20'd0 ) |
 ( (snoop_in == cam_loc709[14:0]) ? cam_loc709 : 20'd0 ) |
 ( (snoop_in == cam_loc710[14:0]) ? cam_loc710 : 20'd0 ) |
 ( (snoop_in == cam_loc711[14:0]) ? cam_loc711 : 20'd0 ) |
 ( (snoop_in == cam_loc712[14:0]) ? cam_loc712 : 20'd0 ) |
 ( (snoop_in == cam_loc713[14:0]) ? cam_loc713 : 20'd0 ) |
 ( (snoop_in == cam_loc714[14:0]) ? cam_loc714 : 20'd0 ) |
 ( (snoop_in == cam_loc715[14:0]) ? cam_loc715 : 20'd0 ) |
 ( (snoop_in == cam_loc716[14:0]) ? cam_loc716 : 20'd0 ) |
 ( (snoop_in == cam_loc717[14:0]) ? cam_loc717 : 20'd0 ) |
 ( (snoop_in == cam_loc718[14:0]) ? cam_loc718 : 20'd0 ) |
 ( (snoop_in == cam_loc719[14:0]) ? cam_loc719 : 20'd0 ) |
 ( (snoop_in == cam_loc720[14:0]) ? cam_loc720 : 20'd0 ) |
 ( (snoop_in == cam_loc721[14:0]) ? cam_loc721 : 20'd0 ) |
 ( (snoop_in == cam_loc722[14:0]) ? cam_loc722 : 20'd0 ) |
 ( (snoop_in == cam_loc723[14:0]) ? cam_loc723 : 20'd0 ) |
 ( (snoop_in == cam_loc724[14:0]) ? cam_loc724 : 20'd0 ) |
 ( (snoop_in == cam_loc725[14:0]) ? cam_loc725 : 20'd0 ) |
 ( (snoop_in == cam_loc726[14:0]) ? cam_loc726 : 20'd0 ) |
 ( (snoop_in == cam_loc727[14:0]) ? cam_loc727 : 20'd0 ) |
 ( (snoop_in == cam_loc728[14:0]) ? cam_loc728 : 20'd0 ) |
 ( (snoop_in == cam_loc729[14:0]) ? cam_loc729 : 20'd0 ) |
 ( (snoop_in == cam_loc730[14:0]) ? cam_loc730 : 20'd0 ) |
 ( (snoop_in == cam_loc731[14:0]) ? cam_loc731 : 20'd0 ) |
 ( (snoop_in == cam_loc732[14:0]) ? cam_loc732 : 20'd0 ) |
 ( (snoop_in == cam_loc733[14:0]) ? cam_loc733 : 20'd0 ) |
 ( (snoop_in == cam_loc734[14:0]) ? cam_loc734 : 20'd0 ) |
 ( (snoop_in == cam_loc735[14:0]) ? cam_loc735 : 20'd0 ) |
 ( (snoop_in == cam_loc736[14:0]) ? cam_loc736 : 20'd0 ) |
 ( (snoop_in == cam_loc737[14:0]) ? cam_loc737 : 20'd0 ) |
 ( (snoop_in == cam_loc738[14:0]) ? cam_loc738 : 20'd0 ) |
 ( (snoop_in == cam_loc739[14:0]) ? cam_loc739 : 20'd0 ) |
 ( (snoop_in == cam_loc740[14:0]) ? cam_loc740 : 20'd0 ) |
 ( (snoop_in == cam_loc741[14:0]) ? cam_loc741 : 20'd0 ) |
 ( (snoop_in == cam_loc742[14:0]) ? cam_loc742 : 20'd0 ) |
 ( (snoop_in == cam_loc743[14:0]) ? cam_loc743 : 20'd0 ) |
 ( (snoop_in == cam_loc744[14:0]) ? cam_loc744 : 20'd0 ) |
 ( (snoop_in == cam_loc745[14:0]) ? cam_loc745 : 20'd0 ) |
 ( (snoop_in == cam_loc746[14:0]) ? cam_loc746 : 20'd0 ) |
 ( (snoop_in == cam_loc747[14:0]) ? cam_loc747 : 20'd0 ) |
 ( (snoop_in == cam_loc748[14:0]) ? cam_loc748 : 20'd0 ) |
 ( (snoop_in == cam_loc749[14:0]) ? cam_loc749 : 20'd0 ) |
 ( (snoop_in == cam_loc750[14:0]) ? cam_loc750 : 20'd0 ) |
 ( (snoop_in == cam_loc751[14:0]) ? cam_loc751 : 20'd0 ) |
 ( (snoop_in == cam_loc752[14:0]) ? cam_loc752 : 20'd0 ) |
 ( (snoop_in == cam_loc753[14:0]) ? cam_loc753 : 20'd0 ) |
 ( (snoop_in == cam_loc754[14:0]) ? cam_loc754 : 20'd0 ) |
 ( (snoop_in == cam_loc755[14:0]) ? cam_loc755 : 20'd0 ) |
 ( (snoop_in == cam_loc756[14:0]) ? cam_loc756 : 20'd0 ) |
 ( (snoop_in == cam_loc757[14:0]) ? cam_loc757 : 20'd0 ) |
 ( (snoop_in == cam_loc758[14:0]) ? cam_loc758 : 20'd0 ) |
 ( (snoop_in == cam_loc759[14:0]) ? cam_loc759 : 20'd0 ) |
 ( (snoop_in == cam_loc760[14:0]) ? cam_loc760 : 20'd0 ) |
 ( (snoop_in == cam_loc761[14:0]) ? cam_loc761 : 20'd0 ) |
 ( (snoop_in == cam_loc762[14:0]) ? cam_loc762 : 20'd0 ) |
 ( (snoop_in == cam_loc763[14:0]) ? cam_loc763 : 20'd0 ) |
 ( (snoop_in == cam_loc764[14:0]) ? cam_loc764 : 20'd0 ) |
 ( (snoop_in == cam_loc765[14:0]) ? cam_loc765 : 20'd0 ) |
 ( (snoop_in == cam_loc766[14:0]) ? cam_loc766 : 20'd0 ) |
 ( (snoop_in == cam_loc767[14:0]) ? cam_loc767 : 20'd0 ) |
 ( (snoop_in == cam_loc768[14:0]) ? cam_loc768 : 20'd0 ) |
 ( (snoop_in == cam_loc769[14:0]) ? cam_loc769 : 20'd0 ) |
 ( (snoop_in == cam_loc770[14:0]) ? cam_loc770 : 20'd0 ) |
 ( (snoop_in == cam_loc771[14:0]) ? cam_loc771 : 20'd0 ) |
 ( (snoop_in == cam_loc772[14:0]) ? cam_loc772 : 20'd0 ) |
 ( (snoop_in == cam_loc773[14:0]) ? cam_loc773 : 20'd0 ) |
 ( (snoop_in == cam_loc774[14:0]) ? cam_loc774 : 20'd0 ) |
 ( (snoop_in == cam_loc775[14:0]) ? cam_loc775 : 20'd0 ) |
 ( (snoop_in == cam_loc776[14:0]) ? cam_loc776 : 20'd0 ) |
 ( (snoop_in == cam_loc777[14:0]) ? cam_loc777 : 20'd0 ) |
 ( (snoop_in == cam_loc778[14:0]) ? cam_loc778 : 20'd0 ) |
 ( (snoop_in == cam_loc779[14:0]) ? cam_loc779 : 20'd0 ) |
 ( (snoop_in == cam_loc780[14:0]) ? cam_loc780 : 20'd0 ) |
 ( (snoop_in == cam_loc781[14:0]) ? cam_loc781 : 20'd0 ) |
 ( (snoop_in == cam_loc782[14:0]) ? cam_loc782 : 20'd0 ) |
 ( (snoop_in == cam_loc783[14:0]) ? cam_loc783 : 20'd0 ) |
 ( (snoop_in == cam_loc784[14:0]) ? cam_loc784 : 20'd0 ) |
 ( (snoop_in == cam_loc785[14:0]) ? cam_loc785 : 20'd0 ) |
 ( (snoop_in == cam_loc786[14:0]) ? cam_loc786 : 20'd0 ) |
 ( (snoop_in == cam_loc787[14:0]) ? cam_loc787 : 20'd0 ) |
 ( (snoop_in == cam_loc788[14:0]) ? cam_loc788 : 20'd0 ) |
 ( (snoop_in == cam_loc789[14:0]) ? cam_loc789 : 20'd0 ) |
 ( (snoop_in == cam_loc790[14:0]) ? cam_loc790 : 20'd0 ) |
 ( (snoop_in == cam_loc791[14:0]) ? cam_loc791 : 20'd0 ) |
 ( (snoop_in == cam_loc792[14:0]) ? cam_loc792 : 20'd0 ) |
 ( (snoop_in == cam_loc793[14:0]) ? cam_loc793 : 20'd0 ) |
 ( (snoop_in == cam_loc794[14:0]) ? cam_loc794 : 20'd0 ) |
 ( (snoop_in == cam_loc795[14:0]) ? cam_loc795 : 20'd0 ) |
 ( (snoop_in == cam_loc796[14:0]) ? cam_loc796 : 20'd0 ) |
 ( (snoop_in == cam_loc797[14:0]) ? cam_loc797 : 20'd0 ) |
 ( (snoop_in == cam_loc798[14:0]) ? cam_loc798 : 20'd0 ) |
 ( (snoop_in == cam_loc799[14:0]) ? cam_loc799 : 20'd0 ) |
 ( (snoop_in == cam_loc800[14:0]) ? cam_loc800 : 20'd0 ) |
 ( (snoop_in == cam_loc801[14:0]) ? cam_loc801 : 20'd0 ) |
 ( (snoop_in == cam_loc802[14:0]) ? cam_loc802 : 20'd0 ) |
 ( (snoop_in == cam_loc803[14:0]) ? cam_loc803 : 20'd0 ) |
 ( (snoop_in == cam_loc804[14:0]) ? cam_loc804 : 20'd0 ) |
 ( (snoop_in == cam_loc805[14:0]) ? cam_loc805 : 20'd0 ) |
 ( (snoop_in == cam_loc806[14:0]) ? cam_loc806 : 20'd0 ) |
 ( (snoop_in == cam_loc807[14:0]) ? cam_loc807 : 20'd0 ) |
 ( (snoop_in == cam_loc808[14:0]) ? cam_loc808 : 20'd0 ) |
 ( (snoop_in == cam_loc809[14:0]) ? cam_loc809 : 20'd0 ) |
 ( (snoop_in == cam_loc810[14:0]) ? cam_loc810 : 20'd0 ) |
 ( (snoop_in == cam_loc811[14:0]) ? cam_loc811 : 20'd0 ) |
 ( (snoop_in == cam_loc812[14:0]) ? cam_loc812 : 20'd0 ) |
 ( (snoop_in == cam_loc813[14:0]) ? cam_loc813 : 20'd0 ) |
 ( (snoop_in == cam_loc814[14:0]) ? cam_loc814 : 20'd0 ) |
 ( (snoop_in == cam_loc815[14:0]) ? cam_loc815 : 20'd0 ) |
 ( (snoop_in == cam_loc816[14:0]) ? cam_loc816 : 20'd0 ) |
 ( (snoop_in == cam_loc817[14:0]) ? cam_loc817 : 20'd0 ) |
 ( (snoop_in == cam_loc818[14:0]) ? cam_loc818 : 20'd0 ) |
 ( (snoop_in == cam_loc819[14:0]) ? cam_loc819 : 20'd0 ) |
 ( (snoop_in == cam_loc820[14:0]) ? cam_loc820 : 20'd0 ) |
 ( (snoop_in == cam_loc821[14:0]) ? cam_loc821 : 20'd0 ) |
 ( (snoop_in == cam_loc822[14:0]) ? cam_loc822 : 20'd0 ) |
 ( (snoop_in == cam_loc823[14:0]) ? cam_loc823 : 20'd0 ) |
 ( (snoop_in == cam_loc824[14:0]) ? cam_loc824 : 20'd0 ) |
 ( (snoop_in == cam_loc825[14:0]) ? cam_loc825 : 20'd0 ) |
 ( (snoop_in == cam_loc826[14:0]) ? cam_loc826 : 20'd0 ) |
 ( (snoop_in == cam_loc827[14:0]) ? cam_loc827 : 20'd0 ) |
 ( (snoop_in == cam_loc828[14:0]) ? cam_loc828 : 20'd0 ) |
 ( (snoop_in == cam_loc829[14:0]) ? cam_loc829 : 20'd0 ) |
 ( (snoop_in == cam_loc830[14:0]) ? cam_loc830 : 20'd0 ) |
 ( (snoop_in == cam_loc831[14:0]) ? cam_loc831 : 20'd0 ) |
 ( (snoop_in == cam_loc832[14:0]) ? cam_loc832 : 20'd0 ) |
 ( (snoop_in == cam_loc833[14:0]) ? cam_loc833 : 20'd0 ) |
 ( (snoop_in == cam_loc834[14:0]) ? cam_loc834 : 20'd0 ) |
 ( (snoop_in == cam_loc835[14:0]) ? cam_loc835 : 20'd0 ) |
 ( (snoop_in == cam_loc836[14:0]) ? cam_loc836 : 20'd0 ) |
 ( (snoop_in == cam_loc837[14:0]) ? cam_loc837 : 20'd0 ) |
 ( (snoop_in == cam_loc838[14:0]) ? cam_loc838 : 20'd0 ) |
 ( (snoop_in == cam_loc839[14:0]) ? cam_loc839 : 20'd0 ) |
 ( (snoop_in == cam_loc840[14:0]) ? cam_loc840 : 20'd0 ) |
 ( (snoop_in == cam_loc841[14:0]) ? cam_loc841 : 20'd0 ) |
 ( (snoop_in == cam_loc842[14:0]) ? cam_loc842 : 20'd0 ) |
 ( (snoop_in == cam_loc843[14:0]) ? cam_loc843 : 20'd0 ) |
 ( (snoop_in == cam_loc844[14:0]) ? cam_loc844 : 20'd0 ) |
 ( (snoop_in == cam_loc845[14:0]) ? cam_loc845 : 20'd0 ) |
 ( (snoop_in == cam_loc846[14:0]) ? cam_loc846 : 20'd0 ) |
 ( (snoop_in == cam_loc847[14:0]) ? cam_loc847 : 20'd0 ) |
 ( (snoop_in == cam_loc848[14:0]) ? cam_loc848 : 20'd0 ) |
 ( (snoop_in == cam_loc849[14:0]) ? cam_loc849 : 20'd0 ) |
 ( (snoop_in == cam_loc850[14:0]) ? cam_loc850 : 20'd0 ) |
 ( (snoop_in == cam_loc851[14:0]) ? cam_loc851 : 20'd0 ) |
 ( (snoop_in == cam_loc852[14:0]) ? cam_loc852 : 20'd0 ) |
 ( (snoop_in == cam_loc853[14:0]) ? cam_loc853 : 20'd0 ) |
 ( (snoop_in == cam_loc854[14:0]) ? cam_loc854 : 20'd0 ) |
 ( (snoop_in == cam_loc855[14:0]) ? cam_loc855 : 20'd0 ) |
 ( (snoop_in == cam_loc856[14:0]) ? cam_loc856 : 20'd0 ) |
 ( (snoop_in == cam_loc857[14:0]) ? cam_loc857 : 20'd0 ) |
 ( (snoop_in == cam_loc858[14:0]) ? cam_loc858 : 20'd0 ) |
 ( (snoop_in == cam_loc859[14:0]) ? cam_loc859 : 20'd0 ) |
 ( (snoop_in == cam_loc860[14:0]) ? cam_loc860 : 20'd0 ) |
 ( (snoop_in == cam_loc861[14:0]) ? cam_loc861 : 20'd0 ) |
 ( (snoop_in == cam_loc862[14:0]) ? cam_loc862 : 20'd0 ) |
 ( (snoop_in == cam_loc863[14:0]) ? cam_loc863 : 20'd0 ) |
 ( (snoop_in == cam_loc864[14:0]) ? cam_loc864 : 20'd0 ) |
 ( (snoop_in == cam_loc865[14:0]) ? cam_loc865 : 20'd0 ) |
 ( (snoop_in == cam_loc866[14:0]) ? cam_loc866 : 20'd0 ) |
 ( (snoop_in == cam_loc867[14:0]) ? cam_loc867 : 20'd0 ) |
 ( (snoop_in == cam_loc868[14:0]) ? cam_loc868 : 20'd0 ) |
 ( (snoop_in == cam_loc869[14:0]) ? cam_loc869 : 20'd0 ) |
 ( (snoop_in == cam_loc870[14:0]) ? cam_loc870 : 20'd0 ) |
 ( (snoop_in == cam_loc871[14:0]) ? cam_loc871 : 20'd0 ) |
 ( (snoop_in == cam_loc872[14:0]) ? cam_loc872 : 20'd0 ) |
 ( (snoop_in == cam_loc873[14:0]) ? cam_loc873 : 20'd0 ) |
 ( (snoop_in == cam_loc874[14:0]) ? cam_loc874 : 20'd0 ) |
 ( (snoop_in == cam_loc875[14:0]) ? cam_loc875 : 20'd0 ) |
 ( (snoop_in == cam_loc876[14:0]) ? cam_loc876 : 20'd0 ) |
 ( (snoop_in == cam_loc877[14:0]) ? cam_loc877 : 20'd0 ) |
 ( (snoop_in == cam_loc878[14:0]) ? cam_loc878 : 20'd0 ) |
 ( (snoop_in == cam_loc879[14:0]) ? cam_loc879 : 20'd0 ) |
 ( (snoop_in == cam_loc880[14:0]) ? cam_loc880 : 20'd0 ) |
 ( (snoop_in == cam_loc881[14:0]) ? cam_loc881 : 20'd0 ) |
 ( (snoop_in == cam_loc882[14:0]) ? cam_loc882 : 20'd0 ) |
 ( (snoop_in == cam_loc883[14:0]) ? cam_loc883 : 20'd0 ) |
 ( (snoop_in == cam_loc884[14:0]) ? cam_loc884 : 20'd0 ) |
 ( (snoop_in == cam_loc885[14:0]) ? cam_loc885 : 20'd0 ) |
 ( (snoop_in == cam_loc886[14:0]) ? cam_loc886 : 20'd0 ) |
 ( (snoop_in == cam_loc887[14:0]) ? cam_loc887 : 20'd0 ) |
 ( (snoop_in == cam_loc888[14:0]) ? cam_loc888 : 20'd0 ) |
 ( (snoop_in == cam_loc889[14:0]) ? cam_loc889 : 20'd0 ) |
 ( (snoop_in == cam_loc890[14:0]) ? cam_loc890 : 20'd0 ) |
 ( (snoop_in == cam_loc891[14:0]) ? cam_loc891 : 20'd0 ) |
 ( (snoop_in == cam_loc892[14:0]) ? cam_loc892 : 20'd0 ) |
 ( (snoop_in == cam_loc893[14:0]) ? cam_loc893 : 20'd0 ) |
 ( (snoop_in == cam_loc894[14:0]) ? cam_loc894 : 20'd0 ) |
 ( (snoop_in == cam_loc895[14:0]) ? cam_loc895 : 20'd0 ) |
 ( (snoop_in == cam_loc896[14:0]) ? cam_loc896 : 20'd0 ) |
 ( (snoop_in == cam_loc897[14:0]) ? cam_loc897 : 20'd0 ) |
 ( (snoop_in == cam_loc898[14:0]) ? cam_loc898 : 20'd0 ) |
 ( (snoop_in == cam_loc899[14:0]) ? cam_loc899 : 20'd0 ) |
 ( (snoop_in == cam_loc900[14:0]) ? cam_loc900 : 20'd0 ) |
 ( (snoop_in == cam_loc901[14:0]) ? cam_loc901 : 20'd0 ) |
 ( (snoop_in == cam_loc902[14:0]) ? cam_loc902 : 20'd0 ) |
 ( (snoop_in == cam_loc903[14:0]) ? cam_loc903 : 20'd0 ) |
 ( (snoop_in == cam_loc904[14:0]) ? cam_loc904 : 20'd0 ) |
 ( (snoop_in == cam_loc905[14:0]) ? cam_loc905 : 20'd0 ) |
 ( (snoop_in == cam_loc906[14:0]) ? cam_loc906 : 20'd0 ) |
 ( (snoop_in == cam_loc907[14:0]) ? cam_loc907 : 20'd0 ) |
 ( (snoop_in == cam_loc908[14:0]) ? cam_loc908 : 20'd0 ) |
 ( (snoop_in == cam_loc909[14:0]) ? cam_loc909 : 20'd0 ) |
 ( (snoop_in == cam_loc910[14:0]) ? cam_loc910 : 20'd0 ) |
 ( (snoop_in == cam_loc911[14:0]) ? cam_loc911 : 20'd0 ) |
 ( (snoop_in == cam_loc912[14:0]) ? cam_loc912 : 20'd0 ) |
 ( (snoop_in == cam_loc913[14:0]) ? cam_loc913 : 20'd0 ) |
 ( (snoop_in == cam_loc914[14:0]) ? cam_loc914 : 20'd0 ) |
 ( (snoop_in == cam_loc915[14:0]) ? cam_loc915 : 20'd0 ) |
 ( (snoop_in == cam_loc916[14:0]) ? cam_loc916 : 20'd0 ) |
 ( (snoop_in == cam_loc917[14:0]) ? cam_loc917 : 20'd0 ) |
 ( (snoop_in == cam_loc918[14:0]) ? cam_loc918 : 20'd0 ) |
 ( (snoop_in == cam_loc919[14:0]) ? cam_loc919 : 20'd0 ) |
 ( (snoop_in == cam_loc920[14:0]) ? cam_loc920 : 20'd0 ) |
 ( (snoop_in == cam_loc921[14:0]) ? cam_loc921 : 20'd0 ) |
 ( (snoop_in == cam_loc922[14:0]) ? cam_loc922 : 20'd0 ) |
 ( (snoop_in == cam_loc923[14:0]) ? cam_loc923 : 20'd0 ) |
 ( (snoop_in == cam_loc924[14:0]) ? cam_loc924 : 20'd0 ) |
 ( (snoop_in == cam_loc925[14:0]) ? cam_loc925 : 20'd0 ) |
 ( (snoop_in == cam_loc926[14:0]) ? cam_loc926 : 20'd0 ) |
 ( (snoop_in == cam_loc927[14:0]) ? cam_loc927 : 20'd0 ) |
 ( (snoop_in == cam_loc928[14:0]) ? cam_loc928 : 20'd0 ) |
 ( (snoop_in == cam_loc929[14:0]) ? cam_loc929 : 20'd0 ) |
 ( (snoop_in == cam_loc930[14:0]) ? cam_loc930 : 20'd0 ) |
 ( (snoop_in == cam_loc931[14:0]) ? cam_loc931 : 20'd0 ) |
 ( (snoop_in == cam_loc932[14:0]) ? cam_loc932 : 20'd0 ) |
 ( (snoop_in == cam_loc933[14:0]) ? cam_loc933 : 20'd0 ) |
 ( (snoop_in == cam_loc934[14:0]) ? cam_loc934 : 20'd0 ) |
 ( (snoop_in == cam_loc935[14:0]) ? cam_loc935 : 20'd0 ) |
 ( (snoop_in == cam_loc936[14:0]) ? cam_loc936 : 20'd0 ) |
 ( (snoop_in == cam_loc937[14:0]) ? cam_loc937 : 20'd0 ) |
 ( (snoop_in == cam_loc938[14:0]) ? cam_loc938 : 20'd0 ) |
 ( (snoop_in == cam_loc939[14:0]) ? cam_loc939 : 20'd0 ) |
 ( (snoop_in == cam_loc940[14:0]) ? cam_loc940 : 20'd0 ) |
 ( (snoop_in == cam_loc941[14:0]) ? cam_loc941 : 20'd0 ) |
 ( (snoop_in == cam_loc942[14:0]) ? cam_loc942 : 20'd0 ) |
 ( (snoop_in == cam_loc943[14:0]) ? cam_loc943 : 20'd0 ) |
 ( (snoop_in == cam_loc944[14:0]) ? cam_loc944 : 20'd0 ) |
 ( (snoop_in == cam_loc945[14:0]) ? cam_loc945 : 20'd0 ) |
 ( (snoop_in == cam_loc946[14:0]) ? cam_loc946 : 20'd0 ) |
 ( (snoop_in == cam_loc947[14:0]) ? cam_loc947 : 20'd0 ) |
 ( (snoop_in == cam_loc948[14:0]) ? cam_loc948 : 20'd0 ) |
 ( (snoop_in == cam_loc949[14:0]) ? cam_loc949 : 20'd0 ) |
 ( (snoop_in == cam_loc950[14:0]) ? cam_loc950 : 20'd0 ) |
 ( (snoop_in == cam_loc951[14:0]) ? cam_loc951 : 20'd0 ) |
 ( (snoop_in == cam_loc952[14:0]) ? cam_loc952 : 20'd0 ) |
 ( (snoop_in == cam_loc953[14:0]) ? cam_loc953 : 20'd0 ) |
 ( (snoop_in == cam_loc954[14:0]) ? cam_loc954 : 20'd0 ) |
 ( (snoop_in == cam_loc955[14:0]) ? cam_loc955 : 20'd0 ) |
 ( (snoop_in == cam_loc956[14:0]) ? cam_loc956 : 20'd0 ) |
 ( (snoop_in == cam_loc957[14:0]) ? cam_loc957 : 20'd0 ) |
 ( (snoop_in == cam_loc958[14:0]) ? cam_loc958 : 20'd0 ) |
 ( (snoop_in == cam_loc959[14:0]) ? cam_loc959 : 20'd0 ) |
 ( (snoop_in == cam_loc960[14:0]) ? cam_loc960 : 20'd0 ) |
 ( (snoop_in == cam_loc961[14:0]) ? cam_loc961 : 20'd0 ) |
 ( (snoop_in == cam_loc962[14:0]) ? cam_loc962 : 20'd0 ) |
 ( (snoop_in == cam_loc963[14:0]) ? cam_loc963 : 20'd0 ) |
 ( (snoop_in == cam_loc964[14:0]) ? cam_loc964 : 20'd0 ) |
 ( (snoop_in == cam_loc965[14:0]) ? cam_loc965 : 20'd0 ) |
 ( (snoop_in == cam_loc966[14:0]) ? cam_loc966 : 20'd0 ) |
 ( (snoop_in == cam_loc967[14:0]) ? cam_loc967 : 20'd0 ) |
 ( (snoop_in == cam_loc968[14:0]) ? cam_loc968 : 20'd0 ) |
 ( (snoop_in == cam_loc969[14:0]) ? cam_loc969 : 20'd0 ) |
 ( (snoop_in == cam_loc970[14:0]) ? cam_loc970 : 20'd0 ) |
 ( (snoop_in == cam_loc971[14:0]) ? cam_loc971 : 20'd0 ) |
 ( (snoop_in == cam_loc972[14:0]) ? cam_loc972 : 20'd0 ) |
 ( (snoop_in == cam_loc973[14:0]) ? cam_loc973 : 20'd0 ) |
 ( (snoop_in == cam_loc974[14:0]) ? cam_loc974 : 20'd0 ) |
 ( (snoop_in == cam_loc975[14:0]) ? cam_loc975 : 20'd0 ) |
 ( (snoop_in == cam_loc976[14:0]) ? cam_loc976 : 20'd0 ) |
 ( (snoop_in == cam_loc977[14:0]) ? cam_loc977 : 20'd0 ) |
 ( (snoop_in == cam_loc978[14:0]) ? cam_loc978 : 20'd0 ) |
 ( (snoop_in == cam_loc979[14:0]) ? cam_loc979 : 20'd0 ) |
 ( (snoop_in == cam_loc980[14:0]) ? cam_loc980 : 20'd0 ) |
 ( (snoop_in == cam_loc981[14:0]) ? cam_loc981 : 20'd0 ) |
 ( (snoop_in == cam_loc982[14:0]) ? cam_loc982 : 20'd0 ) |
 ( (snoop_in == cam_loc983[14:0]) ? cam_loc983 : 20'd0 ) |
 ( (snoop_in == cam_loc984[14:0]) ? cam_loc984 : 20'd0 ) |
 ( (snoop_in == cam_loc985[14:0]) ? cam_loc985 : 20'd0 ) |
 ( (snoop_in == cam_loc986[14:0]) ? cam_loc986 : 20'd0 ) |
 ( (snoop_in == cam_loc987[14:0]) ? cam_loc987 : 20'd0 ) |
 ( (snoop_in == cam_loc988[14:0]) ? cam_loc988 : 20'd0 ) |
 ( (snoop_in == cam_loc989[14:0]) ? cam_loc989 : 20'd0 ) |
 ( (snoop_in == cam_loc990[14:0]) ? cam_loc990 : 20'd0 ) |
 ( (snoop_in == cam_loc991[14:0]) ? cam_loc991 : 20'd0 ) |
 ( (snoop_in == cam_loc992[14:0]) ? cam_loc992 : 20'd0 ) |
 ( (snoop_in == cam_loc993[14:0]) ? cam_loc993 : 20'd0 ) |
 ( (snoop_in == cam_loc994[14:0]) ? cam_loc994 : 20'd0 ) |
 ( (snoop_in == cam_loc995[14:0]) ? cam_loc995 : 20'd0 ) |
 ( (snoop_in == cam_loc996[14:0]) ? cam_loc996 : 20'd0 ) |
 ( (snoop_in == cam_loc997[14:0]) ? cam_loc997 : 20'd0 ) |
 ( (snoop_in == cam_loc998[14:0]) ? cam_loc998 : 20'd0 ) |
 ( (snoop_in == cam_loc999[14:0]) ? cam_loc999 : 20'd0 ) |
 ( (snoop_in == cam_loc1000[14:0]) ? cam_loc1000 : 20'd0 ) |
 ( (snoop_in == cam_loc1001[14:0]) ? cam_loc1001 : 20'd0 ) |
 ( (snoop_in == cam_loc1002[14:0]) ? cam_loc1002 : 20'd0 ) |
 ( (snoop_in == cam_loc1003[14:0]) ? cam_loc1003 : 20'd0 ) |
 ( (snoop_in == cam_loc1004[14:0]) ? cam_loc1004 : 20'd0 ) |
 ( (snoop_in == cam_loc1005[14:0]) ? cam_loc1005 : 20'd0 ) |
 ( (snoop_in == cam_loc1006[14:0]) ? cam_loc1006 : 20'd0 ) |
 ( (snoop_in == cam_loc1007[14:0]) ? cam_loc1007 : 20'd0 ) |
 ( (snoop_in == cam_loc1008[14:0]) ? cam_loc1008 : 20'd0 ) |
 ( (snoop_in == cam_loc1009[14:0]) ? cam_loc1009 : 20'd0 ) |
 ( (snoop_in == cam_loc1010[14:0]) ? cam_loc1010 : 20'd0 ) |
 ( (snoop_in == cam_loc1011[14:0]) ? cam_loc1011 : 20'd0 ) |
 ( (snoop_in == cam_loc1012[14:0]) ? cam_loc1012 : 20'd0 ) |
 ( (snoop_in == cam_loc1013[14:0]) ? cam_loc1013 : 20'd0 ) |
 ( (snoop_in == cam_loc1014[14:0]) ? cam_loc1014 : 20'd0 ) |
 ( (snoop_in == cam_loc1015[14:0]) ? cam_loc1015 : 20'd0 ) |
 ( (snoop_in == cam_loc1016[14:0]) ? cam_loc1016 : 20'd0 ) |
 ( (snoop_in == cam_loc1017[14:0]) ? cam_loc1017 : 20'd0 ) |
 ( (snoop_in == cam_loc1018[14:0]) ? cam_loc1018 : 20'd0 ) |
 ( (snoop_in == cam_loc1019[14:0]) ? cam_loc1019 : 20'd0 ) |
 ( (snoop_in == cam_loc1020[14:0]) ? cam_loc1020 : 20'd0 ) |
 ( (snoop_in == cam_loc1021[14:0]) ? cam_loc1021 : 20'd0 ) |
 ( (snoop_in == cam_loc1022[14:0]) ? cam_loc1022 : 20'd0 ) |
 ( (snoop_in == cam_loc1023[14:0]) ? cam_loc1023 : 20'd0 ) |
 ( (snoop_in == cam_loc1024[14:0]) ? cam_loc1024 : 20'd0 ) |
 ( (snoop_in == cam_loc1025[14:0]) ? cam_loc1025 : 20'd0 ) |
 ( (snoop_in == cam_loc1026[14:0]) ? cam_loc1026 : 20'd0 ) |
 ( (snoop_in == cam_loc1027[14:0]) ? cam_loc1027 : 20'd0 ) |
 ( (snoop_in == cam_loc1028[14:0]) ? cam_loc1028 : 20'd0 ) |
 ( (snoop_in == cam_loc1029[14:0]) ? cam_loc1029 : 20'd0 ) |
 ( (snoop_in == cam_loc1030[14:0]) ? cam_loc1030 : 20'd0 ) |
 ( (snoop_in == cam_loc1031[14:0]) ? cam_loc1031 : 20'd0 ) |
 ( (snoop_in == cam_loc1032[14:0]) ? cam_loc1032 : 20'd0 ) |
 ( (snoop_in == cam_loc1033[14:0]) ? cam_loc1033 : 20'd0 ) |
 ( (snoop_in == cam_loc1034[14:0]) ? cam_loc1034 : 20'd0 ) |
 ( (snoop_in == cam_loc1035[14:0]) ? cam_loc1035 : 20'd0 ) |
 ( (snoop_in == cam_loc1036[14:0]) ? cam_loc1036 : 20'd0 ) |
 ( (snoop_in == cam_loc1037[14:0]) ? cam_loc1037 : 20'd0 ) |
 ( (snoop_in == cam_loc1038[14:0]) ? cam_loc1038 : 20'd0 ) |
 ( (snoop_in == cam_loc1039[14:0]) ? cam_loc1039 : 20'd0 ) |
 ( (snoop_in == cam_loc1040[14:0]) ? cam_loc1040 : 20'd0 ) |
 ( (snoop_in == cam_loc1041[14:0]) ? cam_loc1041 : 20'd0 ) |
 ( (snoop_in == cam_loc1042[14:0]) ? cam_loc1042 : 20'd0 ) |
 ( (snoop_in == cam_loc1043[14:0]) ? cam_loc1043 : 20'd0 ) |
 ( (snoop_in == cam_loc1044[14:0]) ? cam_loc1044 : 20'd0 ) |
 ( (snoop_in == cam_loc1045[14:0]) ? cam_loc1045 : 20'd0 ) |
 ( (snoop_in == cam_loc1046[14:0]) ? cam_loc1046 : 20'd0 ) |
 ( (snoop_in == cam_loc1047[14:0]) ? cam_loc1047 : 20'd0 ) |
 ( (snoop_in == cam_loc1048[14:0]) ? cam_loc1048 : 20'd0 ) |
 ( (snoop_in == cam_loc1049[14:0]) ? cam_loc1049 : 20'd0 ) |
 ( (snoop_in == cam_loc1050[14:0]) ? cam_loc1050 : 20'd0 ) |
 ( (snoop_in == cam_loc1051[14:0]) ? cam_loc1051 : 20'd0 ) |
 ( (snoop_in == cam_loc1052[14:0]) ? cam_loc1052 : 20'd0 ) |
 ( (snoop_in == cam_loc1053[14:0]) ? cam_loc1053 : 20'd0 ) |
 ( (snoop_in == cam_loc1054[14:0]) ? cam_loc1054 : 20'd0 ) |
 ( (snoop_in == cam_loc1055[14:0]) ? cam_loc1055 : 20'd0 ) |
 ( (snoop_in == cam_loc1056[14:0]) ? cam_loc1056 : 20'd0 ) |
 ( (snoop_in == cam_loc1057[14:0]) ? cam_loc1057 : 20'd0 ) |
 ( (snoop_in == cam_loc1058[14:0]) ? cam_loc1058 : 20'd0 ) |
 ( (snoop_in == cam_loc1059[14:0]) ? cam_loc1059 : 20'd0 ) |
 ( (snoop_in == cam_loc1060[14:0]) ? cam_loc1060 : 20'd0 ) |
 ( (snoop_in == cam_loc1061[14:0]) ? cam_loc1061 : 20'd0 ) |
 ( (snoop_in == cam_loc1062[14:0]) ? cam_loc1062 : 20'd0 ) |
 ( (snoop_in == cam_loc1063[14:0]) ? cam_loc1063 : 20'd0 ) |
 ( (snoop_in == cam_loc1064[14:0]) ? cam_loc1064 : 20'd0 ) |
 ( (snoop_in == cam_loc1065[14:0]) ? cam_loc1065 : 20'd0 ) |
 ( (snoop_in == cam_loc1066[14:0]) ? cam_loc1066 : 20'd0 ) |
 ( (snoop_in == cam_loc1067[14:0]) ? cam_loc1067 : 20'd0 ) |
 ( (snoop_in == cam_loc1068[14:0]) ? cam_loc1068 : 20'd0 ) |
 ( (snoop_in == cam_loc1069[14:0]) ? cam_loc1069 : 20'd0 ) |
 ( (snoop_in == cam_loc1070[14:0]) ? cam_loc1070 : 20'd0 ) |
 ( (snoop_in == cam_loc1071[14:0]) ? cam_loc1071 : 20'd0 ) |
 ( (snoop_in == cam_loc1072[14:0]) ? cam_loc1072 : 20'd0 ) |
 ( (snoop_in == cam_loc1073[14:0]) ? cam_loc1073 : 20'd0 ) |
 ( (snoop_in == cam_loc1074[14:0]) ? cam_loc1074 : 20'd0 ) |
 ( (snoop_in == cam_loc1075[14:0]) ? cam_loc1075 : 20'd0 ) |
 ( (snoop_in == cam_loc1076[14:0]) ? cam_loc1076 : 20'd0 ) |
 ( (snoop_in == cam_loc1077[14:0]) ? cam_loc1077 : 20'd0 ) |
 ( (snoop_in == cam_loc1078[14:0]) ? cam_loc1078 : 20'd0 ) |
 ( (snoop_in == cam_loc1079[14:0]) ? cam_loc1079 : 20'd0 ) |
 ( (snoop_in == cam_loc1080[14:0]) ? cam_loc1080 : 20'd0 ) |
 ( (snoop_in == cam_loc1081[14:0]) ? cam_loc1081 : 20'd0 ) |
 ( (snoop_in == cam_loc1082[14:0]) ? cam_loc1082 : 20'd0 ) |
 ( (snoop_in == cam_loc1083[14:0]) ? cam_loc1083 : 20'd0 ) |
 ( (snoop_in == cam_loc1084[14:0]) ? cam_loc1084 : 20'd0 ) |
 ( (snoop_in == cam_loc1085[14:0]) ? cam_loc1085 : 20'd0 ) |
 ( (snoop_in == cam_loc1086[14:0]) ? cam_loc1086 : 20'd0 ) |
 ( (snoop_in == cam_loc1087[14:0]) ? cam_loc1087 : 20'd0 ) |
 ( (snoop_in == cam_loc1088[14:0]) ? cam_loc1088 : 20'd0 ) |
 ( (snoop_in == cam_loc1089[14:0]) ? cam_loc1089 : 20'd0 ) |
 ( (snoop_in == cam_loc1090[14:0]) ? cam_loc1090 : 20'd0 ) |
 ( (snoop_in == cam_loc1091[14:0]) ? cam_loc1091 : 20'd0 ) |
 ( (snoop_in == cam_loc1092[14:0]) ? cam_loc1092 : 20'd0 ) |
 ( (snoop_in == cam_loc1093[14:0]) ? cam_loc1093 : 20'd0 ) |
 ( (snoop_in == cam_loc1094[14:0]) ? cam_loc1094 : 20'd0 ) |
 ( (snoop_in == cam_loc1095[14:0]) ? cam_loc1095 : 20'd0 ) |
 ( (snoop_in == cam_loc1096[14:0]) ? cam_loc1096 : 20'd0 ) |
 ( (snoop_in == cam_loc1097[14:0]) ? cam_loc1097 : 20'd0 ) |
 ( (snoop_in == cam_loc1098[14:0]) ? cam_loc1098 : 20'd0 ) |
 ( (snoop_in == cam_loc1099[14:0]) ? cam_loc1099 : 20'd0 )

;

wire assign freeup_loc = 11'd0 |
( (snoop_in == cam_loc0[14:0]) ? cam_loc0 : 11'd0 ) |
 ( (snoop_in == cam_loc1[14:0]) ? cam_loc1 : 11'd1 ) |
 ( (snoop_in == cam_loc2[14:0]) ? cam_loc2 : 11'd2 ) |
 ( (snoop_in == cam_loc3[14:0]) ? cam_loc3 : 11'd3 ) |
 ( (snoop_in == cam_loc4[14:0]) ? cam_loc4 : 11'd4 ) |
 ( (snoop_in == cam_loc5[14:0]) ? cam_loc5 : 11'd5 ) |
 ( (snoop_in == cam_loc6[14:0]) ? cam_loc6 : 11'd6 ) |
 ( (snoop_in == cam_loc7[14:0]) ? cam_loc7 : 11'd7 ) |
 ( (snoop_in == cam_loc8[14:0]) ? cam_loc8 : 11'd8 ) |
 ( (snoop_in == cam_loc9[14:0]) ? cam_loc9 : 11'd9 ) |
 ( (snoop_in == cam_loc10[14:0]) ? cam_loc10 : 11'd10 ) |
 ( (snoop_in == cam_loc11[14:0]) ? cam_loc11 : 11'd11 ) |
 ( (snoop_in == cam_loc12[14:0]) ? cam_loc12 : 11'd12 ) |
 ( (snoop_in == cam_loc13[14:0]) ? cam_loc13 : 11'd13 ) |
 ( (snoop_in == cam_loc14[14:0]) ? cam_loc14 : 11'd14 ) |
 ( (snoop_in == cam_loc15[14:0]) ? cam_loc15 : 11'd15 ) |
 ( (snoop_in == cam_loc16[14:0]) ? cam_loc16 : 11'd16 ) |
 ( (snoop_in == cam_loc17[14:0]) ? cam_loc17 : 11'd17 ) |
 ( (snoop_in == cam_loc18[14:0]) ? cam_loc18 : 11'd18 ) |
 ( (snoop_in == cam_loc19[14:0]) ? cam_loc19 : 11'd19 ) |
 ( (snoop_in == cam_loc20[14:0]) ? cam_loc20 : 11'd20 ) |
 ( (snoop_in == cam_loc21[14:0]) ? cam_loc21 : 11'd21 ) |
 ( (snoop_in == cam_loc22[14:0]) ? cam_loc22 : 11'd22 ) |
 ( (snoop_in == cam_loc23[14:0]) ? cam_loc23 : 11'd23 ) |
 ( (snoop_in == cam_loc24[14:0]) ? cam_loc24 : 11'd24 ) |
 ( (snoop_in == cam_loc25[14:0]) ? cam_loc25 : 11'd25 ) |
 ( (snoop_in == cam_loc26[14:0]) ? cam_loc26 : 11'd26 ) |
 ( (snoop_in == cam_loc27[14:0]) ? cam_loc27 : 11'd27 ) |
 ( (snoop_in == cam_loc28[14:0]) ? cam_loc28 : 11'd28 ) |
 ( (snoop_in == cam_loc29[14:0]) ? cam_loc29 : 11'd29 ) |
 ( (snoop_in == cam_loc30[14:0]) ? cam_loc30 : 11'd30 ) |
 ( (snoop_in == cam_loc31[14:0]) ? cam_loc31 : 11'd31 ) |
 ( (snoop_in == cam_loc32[14:0]) ? cam_loc32 : 11'd32 ) |
 ( (snoop_in == cam_loc33[14:0]) ? cam_loc33 : 11'd33 ) |
 ( (snoop_in == cam_loc34[14:0]) ? cam_loc34 : 11'd34 ) |
 ( (snoop_in == cam_loc35[14:0]) ? cam_loc35 : 11'd35 ) |
 ( (snoop_in == cam_loc36[14:0]) ? cam_loc36 : 11'd36 ) |
 ( (snoop_in == cam_loc37[14:0]) ? cam_loc37 : 11'd37 ) |
 ( (snoop_in == cam_loc38[14:0]) ? cam_loc38 : 11'd38 ) |
 ( (snoop_in == cam_loc39[14:0]) ? cam_loc39 : 11'd39 ) |
 ( (snoop_in == cam_loc40[14:0]) ? cam_loc40 : 11'd40 ) |
 ( (snoop_in == cam_loc41[14:0]) ? cam_loc41 : 11'd41 ) |
 ( (snoop_in == cam_loc42[14:0]) ? cam_loc42 : 11'd42 ) |
 ( (snoop_in == cam_loc43[14:0]) ? cam_loc43 : 11'd43 ) |
 ( (snoop_in == cam_loc44[14:0]) ? cam_loc44 : 11'd44 ) |
 ( (snoop_in == cam_loc45[14:0]) ? cam_loc45 : 11'd45 ) |
 ( (snoop_in == cam_loc46[14:0]) ? cam_loc46 : 11'd46 ) |
 ( (snoop_in == cam_loc47[14:0]) ? cam_loc47 : 11'd47 ) |
 ( (snoop_in == cam_loc48[14:0]) ? cam_loc48 : 11'd48 ) |
 ( (snoop_in == cam_loc49[14:0]) ? cam_loc49 : 11'd49 ) |
 ( (snoop_in == cam_loc50[14:0]) ? cam_loc50 : 11'd50 ) |
 ( (snoop_in == cam_loc51[14:0]) ? cam_loc51 : 11'd51 ) |
 ( (snoop_in == cam_loc52[14:0]) ? cam_loc52 : 11'd52 ) |
 ( (snoop_in == cam_loc53[14:0]) ? cam_loc53 : 11'd53 ) |
 ( (snoop_in == cam_loc54[14:0]) ? cam_loc54 : 11'd54 ) |
 ( (snoop_in == cam_loc55[14:0]) ? cam_loc55 : 11'd55 ) |
 ( (snoop_in == cam_loc56[14:0]) ? cam_loc56 : 11'd56 ) |
 ( (snoop_in == cam_loc57[14:0]) ? cam_loc57 : 11'd57 ) |
 ( (snoop_in == cam_loc58[14:0]) ? cam_loc58 : 11'd58 ) |
 ( (snoop_in == cam_loc59[14:0]) ? cam_loc59 : 11'd59 ) |
 ( (snoop_in == cam_loc60[14:0]) ? cam_loc60 : 11'd60 ) |
 ( (snoop_in == cam_loc61[14:0]) ? cam_loc61 : 11'd61 ) |
 ( (snoop_in == cam_loc62[14:0]) ? cam_loc62 : 11'd62 ) |
 ( (snoop_in == cam_loc63[14:0]) ? cam_loc63 : 11'd63 ) |
 ( (snoop_in == cam_loc64[14:0]) ? cam_loc64 : 11'd64 ) |
 ( (snoop_in == cam_loc65[14:0]) ? cam_loc65 : 11'd65 ) |
 ( (snoop_in == cam_loc66[14:0]) ? cam_loc66 : 11'd66 ) |
 ( (snoop_in == cam_loc67[14:0]) ? cam_loc67 : 11'd67 ) |
 ( (snoop_in == cam_loc68[14:0]) ? cam_loc68 : 11'd68 ) |
 ( (snoop_in == cam_loc69[14:0]) ? cam_loc69 : 11'd69 ) |
 ( (snoop_in == cam_loc70[14:0]) ? cam_loc70 : 11'd70 ) |
 ( (snoop_in == cam_loc71[14:0]) ? cam_loc71 : 11'd71 ) |
 ( (snoop_in == cam_loc72[14:0]) ? cam_loc72 : 11'd72 ) |
 ( (snoop_in == cam_loc73[14:0]) ? cam_loc73 : 11'd73 ) |
 ( (snoop_in == cam_loc74[14:0]) ? cam_loc74 : 11'd74 ) |
 ( (snoop_in == cam_loc75[14:0]) ? cam_loc75 : 11'd75 ) |
 ( (snoop_in == cam_loc76[14:0]) ? cam_loc76 : 11'd76 ) |
 ( (snoop_in == cam_loc77[14:0]) ? cam_loc77 : 11'd77 ) |
 ( (snoop_in == cam_loc78[14:0]) ? cam_loc78 : 11'd78 ) |
 ( (snoop_in == cam_loc79[14:0]) ? cam_loc79 : 11'd79 ) |
 ( (snoop_in == cam_loc80[14:0]) ? cam_loc80 : 11'd80 ) |
 ( (snoop_in == cam_loc81[14:0]) ? cam_loc81 : 11'd81 ) |
 ( (snoop_in == cam_loc82[14:0]) ? cam_loc82 : 11'd82 ) |
 ( (snoop_in == cam_loc83[14:0]) ? cam_loc83 : 11'd83 ) |
 ( (snoop_in == cam_loc84[14:0]) ? cam_loc84 : 11'd84 ) |
 ( (snoop_in == cam_loc85[14:0]) ? cam_loc85 : 11'd85 ) |
 ( (snoop_in == cam_loc86[14:0]) ? cam_loc86 : 11'd86 ) |
 ( (snoop_in == cam_loc87[14:0]) ? cam_loc87 : 11'd87 ) |
 ( (snoop_in == cam_loc88[14:0]) ? cam_loc88 : 11'd88 ) |
 ( (snoop_in == cam_loc89[14:0]) ? cam_loc89 : 11'd89 ) |
 ( (snoop_in == cam_loc90[14:0]) ? cam_loc90 : 11'd90 ) |
 ( (snoop_in == cam_loc91[14:0]) ? cam_loc91 : 11'd91 ) |
 ( (snoop_in == cam_loc92[14:0]) ? cam_loc92 : 11'd92 ) |
 ( (snoop_in == cam_loc93[14:0]) ? cam_loc93 : 11'd93 ) |
 ( (snoop_in == cam_loc94[14:0]) ? cam_loc94 : 11'd94 ) |
 ( (snoop_in == cam_loc95[14:0]) ? cam_loc95 : 11'd95 ) |
 ( (snoop_in == cam_loc96[14:0]) ? cam_loc96 : 11'd96 ) |
 ( (snoop_in == cam_loc97[14:0]) ? cam_loc97 : 11'd97 ) |
 ( (snoop_in == cam_loc98[14:0]) ? cam_loc98 : 11'd98 ) |
 ( (snoop_in == cam_loc99[14:0]) ? cam_loc99 : 11'd99 ) |
 ( (snoop_in == cam_loc100[14:0]) ? cam_loc100 : 11'd100 ) |
 ( (snoop_in == cam_loc101[14:0]) ? cam_loc101 : 11'd101 ) |
 ( (snoop_in == cam_loc102[14:0]) ? cam_loc102 : 11'd102 ) |
 ( (snoop_in == cam_loc103[14:0]) ? cam_loc103 : 11'd103 ) |
 ( (snoop_in == cam_loc104[14:0]) ? cam_loc104 : 11'd104 ) |
 ( (snoop_in == cam_loc105[14:0]) ? cam_loc105 : 11'd105 ) |
 ( (snoop_in == cam_loc106[14:0]) ? cam_loc106 : 11'd106 ) |
 ( (snoop_in == cam_loc107[14:0]) ? cam_loc107 : 11'd107 ) |
 ( (snoop_in == cam_loc108[14:0]) ? cam_loc108 : 11'd108 ) |
 ( (snoop_in == cam_loc109[14:0]) ? cam_loc109 : 11'd109 ) |
 ( (snoop_in == cam_loc110[14:0]) ? cam_loc110 : 11'd110 ) |
 ( (snoop_in == cam_loc111[14:0]) ? cam_loc111 : 11'd111 ) |
 ( (snoop_in == cam_loc112[14:0]) ? cam_loc112 : 11'd112 ) |
 ( (snoop_in == cam_loc113[14:0]) ? cam_loc113 : 11'd113 ) |
 ( (snoop_in == cam_loc114[14:0]) ? cam_loc114 : 11'd114 ) |
 ( (snoop_in == cam_loc115[14:0]) ? cam_loc115 : 11'd115 ) |
 ( (snoop_in == cam_loc116[14:0]) ? cam_loc116 : 11'd116 ) |
 ( (snoop_in == cam_loc117[14:0]) ? cam_loc117 : 11'd117 ) |
 ( (snoop_in == cam_loc118[14:0]) ? cam_loc118 : 11'd118 ) |
 ( (snoop_in == cam_loc119[14:0]) ? cam_loc119 : 11'd119 ) |
 ( (snoop_in == cam_loc120[14:0]) ? cam_loc120 : 11'd120 ) |
 ( (snoop_in == cam_loc121[14:0]) ? cam_loc121 : 11'd121 ) |
 ( (snoop_in == cam_loc122[14:0]) ? cam_loc122 : 11'd122 ) |
 ( (snoop_in == cam_loc123[14:0]) ? cam_loc123 : 11'd123 ) |
 ( (snoop_in == cam_loc124[14:0]) ? cam_loc124 : 11'd124 ) |
 ( (snoop_in == cam_loc125[14:0]) ? cam_loc125 : 11'd125 ) |
 ( (snoop_in == cam_loc126[14:0]) ? cam_loc126 : 11'd126 ) |
 ( (snoop_in == cam_loc127[14:0]) ? cam_loc127 : 11'd127 ) |
 ( (snoop_in == cam_loc128[14:0]) ? cam_loc128 : 11'd128 ) |
 ( (snoop_in == cam_loc129[14:0]) ? cam_loc129 : 11'd129 ) |
 ( (snoop_in == cam_loc130[14:0]) ? cam_loc130 : 11'd130 ) |
 ( (snoop_in == cam_loc131[14:0]) ? cam_loc131 : 11'd131 ) |
 ( (snoop_in == cam_loc132[14:0]) ? cam_loc132 : 11'd132 ) |
 ( (snoop_in == cam_loc133[14:0]) ? cam_loc133 : 11'd133 ) |
 ( (snoop_in == cam_loc134[14:0]) ? cam_loc134 : 11'd134 ) |
 ( (snoop_in == cam_loc135[14:0]) ? cam_loc135 : 11'd135 ) |
 ( (snoop_in == cam_loc136[14:0]) ? cam_loc136 : 11'd136 ) |
 ( (snoop_in == cam_loc137[14:0]) ? cam_loc137 : 11'd137 ) |
 ( (snoop_in == cam_loc138[14:0]) ? cam_loc138 : 11'd138 ) |
 ( (snoop_in == cam_loc139[14:0]) ? cam_loc139 : 11'd139 ) |
 ( (snoop_in == cam_loc140[14:0]) ? cam_loc140 : 11'd140 ) |
 ( (snoop_in == cam_loc141[14:0]) ? cam_loc141 : 11'd141 ) |
 ( (snoop_in == cam_loc142[14:0]) ? cam_loc142 : 11'd142 ) |
 ( (snoop_in == cam_loc143[14:0]) ? cam_loc143 : 11'd143 ) |
 ( (snoop_in == cam_loc144[14:0]) ? cam_loc144 : 11'd144 ) |
 ( (snoop_in == cam_loc145[14:0]) ? cam_loc145 : 11'd145 ) |
 ( (snoop_in == cam_loc146[14:0]) ? cam_loc146 : 11'd146 ) |
 ( (snoop_in == cam_loc147[14:0]) ? cam_loc147 : 11'd147 ) |
 ( (snoop_in == cam_loc148[14:0]) ? cam_loc148 : 11'd148 ) |
 ( (snoop_in == cam_loc149[14:0]) ? cam_loc149 : 11'd149 ) |
 ( (snoop_in == cam_loc150[14:0]) ? cam_loc150 : 11'd150 ) |
 ( (snoop_in == cam_loc151[14:0]) ? cam_loc151 : 11'd151 ) |
 ( (snoop_in == cam_loc152[14:0]) ? cam_loc152 : 11'd152 ) |
 ( (snoop_in == cam_loc153[14:0]) ? cam_loc153 : 11'd153 ) |
 ( (snoop_in == cam_loc154[14:0]) ? cam_loc154 : 11'd154 ) |
 ( (snoop_in == cam_loc155[14:0]) ? cam_loc155 : 11'd155 ) |
 ( (snoop_in == cam_loc156[14:0]) ? cam_loc156 : 11'd156 ) |
 ( (snoop_in == cam_loc157[14:0]) ? cam_loc157 : 11'd157 ) |
 ( (snoop_in == cam_loc158[14:0]) ? cam_loc158 : 11'd158 ) |
 ( (snoop_in == cam_loc159[14:0]) ? cam_loc159 : 11'd159 ) |
 ( (snoop_in == cam_loc160[14:0]) ? cam_loc160 : 11'd160 ) |
 ( (snoop_in == cam_loc161[14:0]) ? cam_loc161 : 11'd161 ) |
 ( (snoop_in == cam_loc162[14:0]) ? cam_loc162 : 11'd162 ) |
 ( (snoop_in == cam_loc163[14:0]) ? cam_loc163 : 11'd163 ) |
 ( (snoop_in == cam_loc164[14:0]) ? cam_loc164 : 11'd164 ) |
 ( (snoop_in == cam_loc165[14:0]) ? cam_loc165 : 11'd165 ) |
 ( (snoop_in == cam_loc166[14:0]) ? cam_loc166 : 11'd166 ) |
 ( (snoop_in == cam_loc167[14:0]) ? cam_loc167 : 11'd167 ) |
 ( (snoop_in == cam_loc168[14:0]) ? cam_loc168 : 11'd168 ) |
 ( (snoop_in == cam_loc169[14:0]) ? cam_loc169 : 11'd169 ) |
 ( (snoop_in == cam_loc170[14:0]) ? cam_loc170 : 11'd170 ) |
 ( (snoop_in == cam_loc171[14:0]) ? cam_loc171 : 11'd171 ) |
 ( (snoop_in == cam_loc172[14:0]) ? cam_loc172 : 11'd172 ) |
 ( (snoop_in == cam_loc173[14:0]) ? cam_loc173 : 11'd173 ) |
 ( (snoop_in == cam_loc174[14:0]) ? cam_loc174 : 11'd174 ) |
 ( (snoop_in == cam_loc175[14:0]) ? cam_loc175 : 11'd175 ) |
 ( (snoop_in == cam_loc176[14:0]) ? cam_loc176 : 11'd176 ) |
 ( (snoop_in == cam_loc177[14:0]) ? cam_loc177 : 11'd177 ) |
 ( (snoop_in == cam_loc178[14:0]) ? cam_loc178 : 11'd178 ) |
 ( (snoop_in == cam_loc179[14:0]) ? cam_loc179 : 11'd179 ) |
 ( (snoop_in == cam_loc180[14:0]) ? cam_loc180 : 11'd180 ) |
 ( (snoop_in == cam_loc181[14:0]) ? cam_loc181 : 11'd181 ) |
 ( (snoop_in == cam_loc182[14:0]) ? cam_loc182 : 11'd182 ) |
 ( (snoop_in == cam_loc183[14:0]) ? cam_loc183 : 11'd183 ) |
 ( (snoop_in == cam_loc184[14:0]) ? cam_loc184 : 11'd184 ) |
 ( (snoop_in == cam_loc185[14:0]) ? cam_loc185 : 11'd185 ) |
 ( (snoop_in == cam_loc186[14:0]) ? cam_loc186 : 11'd186 ) |
 ( (snoop_in == cam_loc187[14:0]) ? cam_loc187 : 11'd187 ) |
 ( (snoop_in == cam_loc188[14:0]) ? cam_loc188 : 11'd188 ) |
 ( (snoop_in == cam_loc189[14:0]) ? cam_loc189 : 11'd189 ) |
 ( (snoop_in == cam_loc190[14:0]) ? cam_loc190 : 11'd190 ) |
 ( (snoop_in == cam_loc191[14:0]) ? cam_loc191 : 11'd191 ) |
 ( (snoop_in == cam_loc192[14:0]) ? cam_loc192 : 11'd192 ) |
 ( (snoop_in == cam_loc193[14:0]) ? cam_loc193 : 11'd193 ) |
 ( (snoop_in == cam_loc194[14:0]) ? cam_loc194 : 11'd194 ) |
 ( (snoop_in == cam_loc195[14:0]) ? cam_loc195 : 11'd195 ) |
 ( (snoop_in == cam_loc196[14:0]) ? cam_loc196 : 11'd196 ) |
 ( (snoop_in == cam_loc197[14:0]) ? cam_loc197 : 11'd197 ) |
 ( (snoop_in == cam_loc198[14:0]) ? cam_loc198 : 11'd198 ) |
 ( (snoop_in == cam_loc199[14:0]) ? cam_loc199 : 11'd199 ) |
 ( (snoop_in == cam_loc200[14:0]) ? cam_loc200 : 11'd200 ) |
 ( (snoop_in == cam_loc201[14:0]) ? cam_loc201 : 11'd201 ) |
 ( (snoop_in == cam_loc202[14:0]) ? cam_loc202 : 11'd202 ) |
 ( (snoop_in == cam_loc203[14:0]) ? cam_loc203 : 11'd203 ) |
 ( (snoop_in == cam_loc204[14:0]) ? cam_loc204 : 11'd204 ) |
 ( (snoop_in == cam_loc205[14:0]) ? cam_loc205 : 11'd205 ) |
 ( (snoop_in == cam_loc206[14:0]) ? cam_loc206 : 11'd206 ) |
 ( (snoop_in == cam_loc207[14:0]) ? cam_loc207 : 11'd207 ) |
 ( (snoop_in == cam_loc208[14:0]) ? cam_loc208 : 11'd208 ) |
 ( (snoop_in == cam_loc209[14:0]) ? cam_loc209 : 11'd209 ) |
 ( (snoop_in == cam_loc210[14:0]) ? cam_loc210 : 11'd210 ) |
 ( (snoop_in == cam_loc211[14:0]) ? cam_loc211 : 11'd211 ) |
 ( (snoop_in == cam_loc212[14:0]) ? cam_loc212 : 11'd212 ) |
 ( (snoop_in == cam_loc213[14:0]) ? cam_loc213 : 11'd213 ) |
 ( (snoop_in == cam_loc214[14:0]) ? cam_loc214 : 11'd214 ) |
 ( (snoop_in == cam_loc215[14:0]) ? cam_loc215 : 11'd215 ) |
 ( (snoop_in == cam_loc216[14:0]) ? cam_loc216 : 11'd216 ) |
 ( (snoop_in == cam_loc217[14:0]) ? cam_loc217 : 11'd217 ) |
 ( (snoop_in == cam_loc218[14:0]) ? cam_loc218 : 11'd218 ) |
 ( (snoop_in == cam_loc219[14:0]) ? cam_loc219 : 11'd219 ) |
 ( (snoop_in == cam_loc220[14:0]) ? cam_loc220 : 11'd220 ) |
 ( (snoop_in == cam_loc221[14:0]) ? cam_loc221 : 11'd221 ) |
 ( (snoop_in == cam_loc222[14:0]) ? cam_loc222 : 11'd222 ) |
 ( (snoop_in == cam_loc223[14:0]) ? cam_loc223 : 11'd223 ) |
 ( (snoop_in == cam_loc224[14:0]) ? cam_loc224 : 11'd224 ) |
 ( (snoop_in == cam_loc225[14:0]) ? cam_loc225 : 11'd225 ) |
 ( (snoop_in == cam_loc226[14:0]) ? cam_loc226 : 11'd226 ) |
 ( (snoop_in == cam_loc227[14:0]) ? cam_loc227 : 11'd227 ) |
 ( (snoop_in == cam_loc228[14:0]) ? cam_loc228 : 11'd228 ) |
 ( (snoop_in == cam_loc229[14:0]) ? cam_loc229 : 11'd229 ) |
 ( (snoop_in == cam_loc230[14:0]) ? cam_loc230 : 11'd230 ) |
 ( (snoop_in == cam_loc231[14:0]) ? cam_loc231 : 11'd231 ) |
 ( (snoop_in == cam_loc232[14:0]) ? cam_loc232 : 11'd232 ) |
 ( (snoop_in == cam_loc233[14:0]) ? cam_loc233 : 11'd233 ) |
 ( (snoop_in == cam_loc234[14:0]) ? cam_loc234 : 11'd234 ) |
 ( (snoop_in == cam_loc235[14:0]) ? cam_loc235 : 11'd235 ) |
 ( (snoop_in == cam_loc236[14:0]) ? cam_loc236 : 11'd236 ) |
 ( (snoop_in == cam_loc237[14:0]) ? cam_loc237 : 11'd237 ) |
 ( (snoop_in == cam_loc238[14:0]) ? cam_loc238 : 11'd238 ) |
 ( (snoop_in == cam_loc239[14:0]) ? cam_loc239 : 11'd239 ) |
 ( (snoop_in == cam_loc240[14:0]) ? cam_loc240 : 11'd240 ) |
 ( (snoop_in == cam_loc241[14:0]) ? cam_loc241 : 11'd241 ) |
 ( (snoop_in == cam_loc242[14:0]) ? cam_loc242 : 11'd242 ) |
 ( (snoop_in == cam_loc243[14:0]) ? cam_loc243 : 11'd243 ) |
 ( (snoop_in == cam_loc244[14:0]) ? cam_loc244 : 11'd244 ) |
 ( (snoop_in == cam_loc245[14:0]) ? cam_loc245 : 11'd245 ) |
 ( (snoop_in == cam_loc246[14:0]) ? cam_loc246 : 11'd246 ) |
 ( (snoop_in == cam_loc247[14:0]) ? cam_loc247 : 11'd247 ) |
 ( (snoop_in == cam_loc248[14:0]) ? cam_loc248 : 11'd248 ) |
 ( (snoop_in == cam_loc249[14:0]) ? cam_loc249 : 11'd249 ) |
 ( (snoop_in == cam_loc250[14:0]) ? cam_loc250 : 11'd250 ) |
 ( (snoop_in == cam_loc251[14:0]) ? cam_loc251 : 11'd251 ) |
 ( (snoop_in == cam_loc252[14:0]) ? cam_loc252 : 11'd252 ) |
 ( (snoop_in == cam_loc253[14:0]) ? cam_loc253 : 11'd253 ) |
 ( (snoop_in == cam_loc254[14:0]) ? cam_loc254 : 11'd254 ) |
 ( (snoop_in == cam_loc255[14:0]) ? cam_loc255 : 11'd255 ) |
 ( (snoop_in == cam_loc256[14:0]) ? cam_loc256 : 11'd256 ) |
 ( (snoop_in == cam_loc257[14:0]) ? cam_loc257 : 11'd257 ) |
 ( (snoop_in == cam_loc258[14:0]) ? cam_loc258 : 11'd258 ) |
 ( (snoop_in == cam_loc259[14:0]) ? cam_loc259 : 11'd259 ) |
 ( (snoop_in == cam_loc260[14:0]) ? cam_loc260 : 11'd260 ) |
 ( (snoop_in == cam_loc261[14:0]) ? cam_loc261 : 11'd261 ) |
 ( (snoop_in == cam_loc262[14:0]) ? cam_loc262 : 11'd262 ) |
 ( (snoop_in == cam_loc263[14:0]) ? cam_loc263 : 11'd263 ) |
 ( (snoop_in == cam_loc264[14:0]) ? cam_loc264 : 11'd264 ) |
 ( (snoop_in == cam_loc265[14:0]) ? cam_loc265 : 11'd265 ) |
 ( (snoop_in == cam_loc266[14:0]) ? cam_loc266 : 11'd266 ) |
 ( (snoop_in == cam_loc267[14:0]) ? cam_loc267 : 11'd267 ) |
 ( (snoop_in == cam_loc268[14:0]) ? cam_loc268 : 11'd268 ) |
 ( (snoop_in == cam_loc269[14:0]) ? cam_loc269 : 11'd269 ) |
 ( (snoop_in == cam_loc270[14:0]) ? cam_loc270 : 11'd270 ) |
 ( (snoop_in == cam_loc271[14:0]) ? cam_loc271 : 11'd271 ) |
 ( (snoop_in == cam_loc272[14:0]) ? cam_loc272 : 11'd272 ) |
 ( (snoop_in == cam_loc273[14:0]) ? cam_loc273 : 11'd273 ) |
 ( (snoop_in == cam_loc274[14:0]) ? cam_loc274 : 11'd274 ) |
 ( (snoop_in == cam_loc275[14:0]) ? cam_loc275 : 11'd275 ) |
 ( (snoop_in == cam_loc276[14:0]) ? cam_loc276 : 11'd276 ) |
 ( (snoop_in == cam_loc277[14:0]) ? cam_loc277 : 11'd277 ) |
 ( (snoop_in == cam_loc278[14:0]) ? cam_loc278 : 11'd278 ) |
 ( (snoop_in == cam_loc279[14:0]) ? cam_loc279 : 11'd279 ) |
 ( (snoop_in == cam_loc280[14:0]) ? cam_loc280 : 11'd280 ) |
 ( (snoop_in == cam_loc281[14:0]) ? cam_loc281 : 11'd281 ) |
 ( (snoop_in == cam_loc282[14:0]) ? cam_loc282 : 11'd282 ) |
 ( (snoop_in == cam_loc283[14:0]) ? cam_loc283 : 11'd283 ) |
 ( (snoop_in == cam_loc284[14:0]) ? cam_loc284 : 11'd284 ) |
 ( (snoop_in == cam_loc285[14:0]) ? cam_loc285 : 11'd285 ) |
 ( (snoop_in == cam_loc286[14:0]) ? cam_loc286 : 11'd286 ) |
 ( (snoop_in == cam_loc287[14:0]) ? cam_loc287 : 11'd287 ) |
 ( (snoop_in == cam_loc288[14:0]) ? cam_loc288 : 11'd288 ) |
 ( (snoop_in == cam_loc289[14:0]) ? cam_loc289 : 11'd289 ) |
 ( (snoop_in == cam_loc290[14:0]) ? cam_loc290 : 11'd290 ) |
 ( (snoop_in == cam_loc291[14:0]) ? cam_loc291 : 11'd291 ) |
 ( (snoop_in == cam_loc292[14:0]) ? cam_loc292 : 11'd292 ) |
 ( (snoop_in == cam_loc293[14:0]) ? cam_loc293 : 11'd293 ) |
 ( (snoop_in == cam_loc294[14:0]) ? cam_loc294 : 11'd294 ) |
 ( (snoop_in == cam_loc295[14:0]) ? cam_loc295 : 11'd295 ) |
 ( (snoop_in == cam_loc296[14:0]) ? cam_loc296 : 11'd296 ) |
 ( (snoop_in == cam_loc297[14:0]) ? cam_loc297 : 11'd297 ) |
 ( (snoop_in == cam_loc298[14:0]) ? cam_loc298 : 11'd298 ) |
 ( (snoop_in == cam_loc299[14:0]) ? cam_loc299 : 11'd299 ) |
 ( (snoop_in == cam_loc300[14:0]) ? cam_loc300 : 11'd300 ) |
 ( (snoop_in == cam_loc301[14:0]) ? cam_loc301 : 11'd301 ) |
 ( (snoop_in == cam_loc302[14:0]) ? cam_loc302 : 11'd302 ) |
 ( (snoop_in == cam_loc303[14:0]) ? cam_loc303 : 11'd303 ) |
 ( (snoop_in == cam_loc304[14:0]) ? cam_loc304 : 11'd304 ) |
 ( (snoop_in == cam_loc305[14:0]) ? cam_loc305 : 11'd305 ) |
 ( (snoop_in == cam_loc306[14:0]) ? cam_loc306 : 11'd306 ) |
 ( (snoop_in == cam_loc307[14:0]) ? cam_loc307 : 11'd307 ) |
 ( (snoop_in == cam_loc308[14:0]) ? cam_loc308 : 11'd308 ) |
 ( (snoop_in == cam_loc309[14:0]) ? cam_loc309 : 11'd309 ) |
 ( (snoop_in == cam_loc310[14:0]) ? cam_loc310 : 11'd310 ) |
 ( (snoop_in == cam_loc311[14:0]) ? cam_loc311 : 11'd311 ) |
 ( (snoop_in == cam_loc312[14:0]) ? cam_loc312 : 11'd312 ) |
 ( (snoop_in == cam_loc313[14:0]) ? cam_loc313 : 11'd313 ) |
 ( (snoop_in == cam_loc314[14:0]) ? cam_loc314 : 11'd314 ) |
 ( (snoop_in == cam_loc315[14:0]) ? cam_loc315 : 11'd315 ) |
 ( (snoop_in == cam_loc316[14:0]) ? cam_loc316 : 11'd316 ) |
 ( (snoop_in == cam_loc317[14:0]) ? cam_loc317 : 11'd317 ) |
 ( (snoop_in == cam_loc318[14:0]) ? cam_loc318 : 11'd318 ) |
 ( (snoop_in == cam_loc319[14:0]) ? cam_loc319 : 11'd319 ) |
 ( (snoop_in == cam_loc320[14:0]) ? cam_loc320 : 11'd320 ) |
 ( (snoop_in == cam_loc321[14:0]) ? cam_loc321 : 11'd321 ) |
 ( (snoop_in == cam_loc322[14:0]) ? cam_loc322 : 11'd322 ) |
 ( (snoop_in == cam_loc323[14:0]) ? cam_loc323 : 11'd323 ) |
 ( (snoop_in == cam_loc324[14:0]) ? cam_loc324 : 11'd324 ) |
 ( (snoop_in == cam_loc325[14:0]) ? cam_loc325 : 11'd325 ) |
 ( (snoop_in == cam_loc326[14:0]) ? cam_loc326 : 11'd326 ) |
 ( (snoop_in == cam_loc327[14:0]) ? cam_loc327 : 11'd327 ) |
 ( (snoop_in == cam_loc328[14:0]) ? cam_loc328 : 11'd328 ) |
 ( (snoop_in == cam_loc329[14:0]) ? cam_loc329 : 11'd329 ) |
 ( (snoop_in == cam_loc330[14:0]) ? cam_loc330 : 11'd330 ) |
 ( (snoop_in == cam_loc331[14:0]) ? cam_loc331 : 11'd331 ) |
 ( (snoop_in == cam_loc332[14:0]) ? cam_loc332 : 11'd332 ) |
 ( (snoop_in == cam_loc333[14:0]) ? cam_loc333 : 11'd333 ) |
 ( (snoop_in == cam_loc334[14:0]) ? cam_loc334 : 11'd334 ) |
 ( (snoop_in == cam_loc335[14:0]) ? cam_loc335 : 11'd335 ) |
 ( (snoop_in == cam_loc336[14:0]) ? cam_loc336 : 11'd336 ) |
 ( (snoop_in == cam_loc337[14:0]) ? cam_loc337 : 11'd337 ) |
 ( (snoop_in == cam_loc338[14:0]) ? cam_loc338 : 11'd338 ) |
 ( (snoop_in == cam_loc339[14:0]) ? cam_loc339 : 11'd339 ) |
 ( (snoop_in == cam_loc340[14:0]) ? cam_loc340 : 11'd340 ) |
 ( (snoop_in == cam_loc341[14:0]) ? cam_loc341 : 11'd341 ) |
 ( (snoop_in == cam_loc342[14:0]) ? cam_loc342 : 11'd342 ) |
 ( (snoop_in == cam_loc343[14:0]) ? cam_loc343 : 11'd343 ) |
 ( (snoop_in == cam_loc344[14:0]) ? cam_loc344 : 11'd344 ) |
 ( (snoop_in == cam_loc345[14:0]) ? cam_loc345 : 11'd345 ) |
 ( (snoop_in == cam_loc346[14:0]) ? cam_loc346 : 11'd346 ) |
 ( (snoop_in == cam_loc347[14:0]) ? cam_loc347 : 11'd347 ) |
 ( (snoop_in == cam_loc348[14:0]) ? cam_loc348 : 11'd348 ) |
 ( (snoop_in == cam_loc349[14:0]) ? cam_loc349 : 11'd349 ) |
 ( (snoop_in == cam_loc350[14:0]) ? cam_loc350 : 11'd350 ) |
 ( (snoop_in == cam_loc351[14:0]) ? cam_loc351 : 11'd351 ) |
 ( (snoop_in == cam_loc352[14:0]) ? cam_loc352 : 11'd352 ) |
 ( (snoop_in == cam_loc353[14:0]) ? cam_loc353 : 11'd353 ) |
 ( (snoop_in == cam_loc354[14:0]) ? cam_loc354 : 11'd354 ) |
 ( (snoop_in == cam_loc355[14:0]) ? cam_loc355 : 11'd355 ) |
 ( (snoop_in == cam_loc356[14:0]) ? cam_loc356 : 11'd356 ) |
 ( (snoop_in == cam_loc357[14:0]) ? cam_loc357 : 11'd357 ) |
 ( (snoop_in == cam_loc358[14:0]) ? cam_loc358 : 11'd358 ) |
 ( (snoop_in == cam_loc359[14:0]) ? cam_loc359 : 11'd359 ) |
 ( (snoop_in == cam_loc360[14:0]) ? cam_loc360 : 11'd360 ) |
 ( (snoop_in == cam_loc361[14:0]) ? cam_loc361 : 11'd361 ) |
 ( (snoop_in == cam_loc362[14:0]) ? cam_loc362 : 11'd362 ) |
 ( (snoop_in == cam_loc363[14:0]) ? cam_loc363 : 11'd363 ) |
 ( (snoop_in == cam_loc364[14:0]) ? cam_loc364 : 11'd364 ) |
 ( (snoop_in == cam_loc365[14:0]) ? cam_loc365 : 11'd365 ) |
 ( (snoop_in == cam_loc366[14:0]) ? cam_loc366 : 11'd366 ) |
 ( (snoop_in == cam_loc367[14:0]) ? cam_loc367 : 11'd367 ) |
 ( (snoop_in == cam_loc368[14:0]) ? cam_loc368 : 11'd368 ) |
 ( (snoop_in == cam_loc369[14:0]) ? cam_loc369 : 11'd369 ) |
 ( (snoop_in == cam_loc370[14:0]) ? cam_loc370 : 11'd370 ) |
 ( (snoop_in == cam_loc371[14:0]) ? cam_loc371 : 11'd371 ) |
 ( (snoop_in == cam_loc372[14:0]) ? cam_loc372 : 11'd372 ) |
 ( (snoop_in == cam_loc373[14:0]) ? cam_loc373 : 11'd373 ) |
 ( (snoop_in == cam_loc374[14:0]) ? cam_loc374 : 11'd374 ) |
 ( (snoop_in == cam_loc375[14:0]) ? cam_loc375 : 11'd375 ) |
 ( (snoop_in == cam_loc376[14:0]) ? cam_loc376 : 11'd376 ) |
 ( (snoop_in == cam_loc377[14:0]) ? cam_loc377 : 11'd377 ) |
 ( (snoop_in == cam_loc378[14:0]) ? cam_loc378 : 11'd378 ) |
 ( (snoop_in == cam_loc379[14:0]) ? cam_loc379 : 11'd379 ) |
 ( (snoop_in == cam_loc380[14:0]) ? cam_loc380 : 11'd380 ) |
 ( (snoop_in == cam_loc381[14:0]) ? cam_loc381 : 11'd381 ) |
 ( (snoop_in == cam_loc382[14:0]) ? cam_loc382 : 11'd382 ) |
 ( (snoop_in == cam_loc383[14:0]) ? cam_loc383 : 11'd383 ) |
 ( (snoop_in == cam_loc384[14:0]) ? cam_loc384 : 11'd384 ) |
 ( (snoop_in == cam_loc385[14:0]) ? cam_loc385 : 11'd385 ) |
 ( (snoop_in == cam_loc386[14:0]) ? cam_loc386 : 11'd386 ) |
 ( (snoop_in == cam_loc387[14:0]) ? cam_loc387 : 11'd387 ) |
 ( (snoop_in == cam_loc388[14:0]) ? cam_loc388 : 11'd388 ) |
 ( (snoop_in == cam_loc389[14:0]) ? cam_loc389 : 11'd389 ) |
 ( (snoop_in == cam_loc390[14:0]) ? cam_loc390 : 11'd390 ) |
 ( (snoop_in == cam_loc391[14:0]) ? cam_loc391 : 11'd391 ) |
 ( (snoop_in == cam_loc392[14:0]) ? cam_loc392 : 11'd392 ) |
 ( (snoop_in == cam_loc393[14:0]) ? cam_loc393 : 11'd393 ) |
 ( (snoop_in == cam_loc394[14:0]) ? cam_loc394 : 11'd394 ) |
 ( (snoop_in == cam_loc395[14:0]) ? cam_loc395 : 11'd395 ) |
 ( (snoop_in == cam_loc396[14:0]) ? cam_loc396 : 11'd396 ) |
 ( (snoop_in == cam_loc397[14:0]) ? cam_loc397 : 11'd397 ) |
 ( (snoop_in == cam_loc398[14:0]) ? cam_loc398 : 11'd398 ) |
 ( (snoop_in == cam_loc399[14:0]) ? cam_loc399 : 11'd399 ) |
 ( (snoop_in == cam_loc400[14:0]) ? cam_loc400 : 11'd400 ) |
 ( (snoop_in == cam_loc401[14:0]) ? cam_loc401 : 11'd401 ) |
 ( (snoop_in == cam_loc402[14:0]) ? cam_loc402 : 11'd402 ) |
 ( (snoop_in == cam_loc403[14:0]) ? cam_loc403 : 11'd403 ) |
 ( (snoop_in == cam_loc404[14:0]) ? cam_loc404 : 11'd404 ) |
 ( (snoop_in == cam_loc405[14:0]) ? cam_loc405 : 11'd405 ) |
 ( (snoop_in == cam_loc406[14:0]) ? cam_loc406 : 11'd406 ) |
 ( (snoop_in == cam_loc407[14:0]) ? cam_loc407 : 11'd407 ) |
 ( (snoop_in == cam_loc408[14:0]) ? cam_loc408 : 11'd408 ) |
 ( (snoop_in == cam_loc409[14:0]) ? cam_loc409 : 11'd409 ) |
 ( (snoop_in == cam_loc410[14:0]) ? cam_loc410 : 11'd410 ) |
 ( (snoop_in == cam_loc411[14:0]) ? cam_loc411 : 11'd411 ) |
 ( (snoop_in == cam_loc412[14:0]) ? cam_loc412 : 11'd412 ) |
 ( (snoop_in == cam_loc413[14:0]) ? cam_loc413 : 11'd413 ) |
 ( (snoop_in == cam_loc414[14:0]) ? cam_loc414 : 11'd414 ) |
 ( (snoop_in == cam_loc415[14:0]) ? cam_loc415 : 11'd415 ) |
 ( (snoop_in == cam_loc416[14:0]) ? cam_loc416 : 11'd416 ) |
 ( (snoop_in == cam_loc417[14:0]) ? cam_loc417 : 11'd417 ) |
 ( (snoop_in == cam_loc418[14:0]) ? cam_loc418 : 11'd418 ) |
 ( (snoop_in == cam_loc419[14:0]) ? cam_loc419 : 11'd419 ) |
 ( (snoop_in == cam_loc420[14:0]) ? cam_loc420 : 11'd420 ) |
 ( (snoop_in == cam_loc421[14:0]) ? cam_loc421 : 11'd421 ) |
 ( (snoop_in == cam_loc422[14:0]) ? cam_loc422 : 11'd422 ) |
 ( (snoop_in == cam_loc423[14:0]) ? cam_loc423 : 11'd423 ) |
 ( (snoop_in == cam_loc424[14:0]) ? cam_loc424 : 11'd424 ) |
 ( (snoop_in == cam_loc425[14:0]) ? cam_loc425 : 11'd425 ) |
 ( (snoop_in == cam_loc426[14:0]) ? cam_loc426 : 11'd426 ) |
 ( (snoop_in == cam_loc427[14:0]) ? cam_loc427 : 11'd427 ) |
 ( (snoop_in == cam_loc428[14:0]) ? cam_loc428 : 11'd428 ) |
 ( (snoop_in == cam_loc429[14:0]) ? cam_loc429 : 11'd429 ) |
 ( (snoop_in == cam_loc430[14:0]) ? cam_loc430 : 11'd430 ) |
 ( (snoop_in == cam_loc431[14:0]) ? cam_loc431 : 11'd431 ) |
 ( (snoop_in == cam_loc432[14:0]) ? cam_loc432 : 11'd432 ) |
 ( (snoop_in == cam_loc433[14:0]) ? cam_loc433 : 11'd433 ) |
 ( (snoop_in == cam_loc434[14:0]) ? cam_loc434 : 11'd434 ) |
 ( (snoop_in == cam_loc435[14:0]) ? cam_loc435 : 11'd435 ) |
 ( (snoop_in == cam_loc436[14:0]) ? cam_loc436 : 11'd436 ) |
 ( (snoop_in == cam_loc437[14:0]) ? cam_loc437 : 11'd437 ) |
 ( (snoop_in == cam_loc438[14:0]) ? cam_loc438 : 11'd438 ) |
 ( (snoop_in == cam_loc439[14:0]) ? cam_loc439 : 11'd439 ) |
 ( (snoop_in == cam_loc440[14:0]) ? cam_loc440 : 11'd440 ) |
 ( (snoop_in == cam_loc441[14:0]) ? cam_loc441 : 11'd441 ) |
 ( (snoop_in == cam_loc442[14:0]) ? cam_loc442 : 11'd442 ) |
 ( (snoop_in == cam_loc443[14:0]) ? cam_loc443 : 11'd443 ) |
 ( (snoop_in == cam_loc444[14:0]) ? cam_loc444 : 11'd444 ) |
 ( (snoop_in == cam_loc445[14:0]) ? cam_loc445 : 11'd445 ) |
 ( (snoop_in == cam_loc446[14:0]) ? cam_loc446 : 11'd446 ) |
 ( (snoop_in == cam_loc447[14:0]) ? cam_loc447 : 11'd447 ) |
 ( (snoop_in == cam_loc448[14:0]) ? cam_loc448 : 11'd448 ) |
 ( (snoop_in == cam_loc449[14:0]) ? cam_loc449 : 11'd449 ) |
 ( (snoop_in == cam_loc450[14:0]) ? cam_loc450 : 11'd450 ) |
 ( (snoop_in == cam_loc451[14:0]) ? cam_loc451 : 11'd451 ) |
 ( (snoop_in == cam_loc452[14:0]) ? cam_loc452 : 11'd452 ) |
 ( (snoop_in == cam_loc453[14:0]) ? cam_loc453 : 11'd453 ) |
 ( (snoop_in == cam_loc454[14:0]) ? cam_loc454 : 11'd454 ) |
 ( (snoop_in == cam_loc455[14:0]) ? cam_loc455 : 11'd455 ) |
 ( (snoop_in == cam_loc456[14:0]) ? cam_loc456 : 11'd456 ) |
 ( (snoop_in == cam_loc457[14:0]) ? cam_loc457 : 11'd457 ) |
 ( (snoop_in == cam_loc458[14:0]) ? cam_loc458 : 11'd458 ) |
 ( (snoop_in == cam_loc459[14:0]) ? cam_loc459 : 11'd459 ) |
 ( (snoop_in == cam_loc460[14:0]) ? cam_loc460 : 11'd460 ) |
 ( (snoop_in == cam_loc461[14:0]) ? cam_loc461 : 11'd461 ) |
 ( (snoop_in == cam_loc462[14:0]) ? cam_loc462 : 11'd462 ) |
 ( (snoop_in == cam_loc463[14:0]) ? cam_loc463 : 11'd463 ) |
 ( (snoop_in == cam_loc464[14:0]) ? cam_loc464 : 11'd464 ) |
 ( (snoop_in == cam_loc465[14:0]) ? cam_loc465 : 11'd465 ) |
 ( (snoop_in == cam_loc466[14:0]) ? cam_loc466 : 11'd466 ) |
 ( (snoop_in == cam_loc467[14:0]) ? cam_loc467 : 11'd467 ) |
 ( (snoop_in == cam_loc468[14:0]) ? cam_loc468 : 11'd468 ) |
 ( (snoop_in == cam_loc469[14:0]) ? cam_loc469 : 11'd469 ) |
 ( (snoop_in == cam_loc470[14:0]) ? cam_loc470 : 11'd470 ) |
 ( (snoop_in == cam_loc471[14:0]) ? cam_loc471 : 11'd471 ) |
 ( (snoop_in == cam_loc472[14:0]) ? cam_loc472 : 11'd472 ) |
 ( (snoop_in == cam_loc473[14:0]) ? cam_loc473 : 11'd473 ) |
 ( (snoop_in == cam_loc474[14:0]) ? cam_loc474 : 11'd474 ) |
 ( (snoop_in == cam_loc475[14:0]) ? cam_loc475 : 11'd475 ) |
 ( (snoop_in == cam_loc476[14:0]) ? cam_loc476 : 11'd476 ) |
 ( (snoop_in == cam_loc477[14:0]) ? cam_loc477 : 11'd477 ) |
 ( (snoop_in == cam_loc478[14:0]) ? cam_loc478 : 11'd478 ) |
 ( (snoop_in == cam_loc479[14:0]) ? cam_loc479 : 11'd479 ) |
 ( (snoop_in == cam_loc480[14:0]) ? cam_loc480 : 11'd480 ) |
 ( (snoop_in == cam_loc481[14:0]) ? cam_loc481 : 11'd481 ) |
 ( (snoop_in == cam_loc482[14:0]) ? cam_loc482 : 11'd482 ) |
 ( (snoop_in == cam_loc483[14:0]) ? cam_loc483 : 11'd483 ) |
 ( (snoop_in == cam_loc484[14:0]) ? cam_loc484 : 11'd484 ) |
 ( (snoop_in == cam_loc485[14:0]) ? cam_loc485 : 11'd485 ) |
 ( (snoop_in == cam_loc486[14:0]) ? cam_loc486 : 11'd486 ) |
 ( (snoop_in == cam_loc487[14:0]) ? cam_loc487 : 11'd487 ) |
 ( (snoop_in == cam_loc488[14:0]) ? cam_loc488 : 11'd488 ) |
 ( (snoop_in == cam_loc489[14:0]) ? cam_loc489 : 11'd489 ) |
 ( (snoop_in == cam_loc490[14:0]) ? cam_loc490 : 11'd490 ) |
 ( (snoop_in == cam_loc491[14:0]) ? cam_loc491 : 11'd491 ) |
 ( (snoop_in == cam_loc492[14:0]) ? cam_loc492 : 11'd492 ) |
 ( (snoop_in == cam_loc493[14:0]) ? cam_loc493 : 11'd493 ) |
 ( (snoop_in == cam_loc494[14:0]) ? cam_loc494 : 11'd494 ) |
 ( (snoop_in == cam_loc495[14:0]) ? cam_loc495 : 11'd495 ) |
 ( (snoop_in == cam_loc496[14:0]) ? cam_loc496 : 11'd496 ) |
 ( (snoop_in == cam_loc497[14:0]) ? cam_loc497 : 11'd497 ) |
 ( (snoop_in == cam_loc498[14:0]) ? cam_loc498 : 11'd498 ) |
 ( (snoop_in == cam_loc499[14:0]) ? cam_loc499 : 11'd499 ) |
 ( (snoop_in == cam_loc500[14:0]) ? cam_loc500 : 11'd500 ) |
 ( (snoop_in == cam_loc501[14:0]) ? cam_loc501 : 11'd501 ) |
 ( (snoop_in == cam_loc502[14:0]) ? cam_loc502 : 11'd502 ) |
 ( (snoop_in == cam_loc503[14:0]) ? cam_loc503 : 11'd503 ) |
 ( (snoop_in == cam_loc504[14:0]) ? cam_loc504 : 11'd504 ) |
 ( (snoop_in == cam_loc505[14:0]) ? cam_loc505 : 11'd505 ) |
 ( (snoop_in == cam_loc506[14:0]) ? cam_loc506 : 11'd506 ) |
 ( (snoop_in == cam_loc507[14:0]) ? cam_loc507 : 11'd507 ) |
 ( (snoop_in == cam_loc508[14:0]) ? cam_loc508 : 11'd508 ) |
 ( (snoop_in == cam_loc509[14:0]) ? cam_loc509 : 11'd509 ) |
 ( (snoop_in == cam_loc510[14:0]) ? cam_loc510 : 11'd510 ) |
 ( (snoop_in == cam_loc511[14:0]) ? cam_loc511 : 11'd511 ) |
 ( (snoop_in == cam_loc512[14:0]) ? cam_loc512 : 11'd512 ) |
 ( (snoop_in == cam_loc513[14:0]) ? cam_loc513 : 11'd513 ) |
 ( (snoop_in == cam_loc514[14:0]) ? cam_loc514 : 11'd514 ) |
 ( (snoop_in == cam_loc515[14:0]) ? cam_loc515 : 11'd515 ) |
 ( (snoop_in == cam_loc516[14:0]) ? cam_loc516 : 11'd516 ) |
 ( (snoop_in == cam_loc517[14:0]) ? cam_loc517 : 11'd517 ) |
 ( (snoop_in == cam_loc518[14:0]) ? cam_loc518 : 11'd518 ) |
 ( (snoop_in == cam_loc519[14:0]) ? cam_loc519 : 11'd519 ) |
 ( (snoop_in == cam_loc520[14:0]) ? cam_loc520 : 11'd520 ) |
 ( (snoop_in == cam_loc521[14:0]) ? cam_loc521 : 11'd521 ) |
 ( (snoop_in == cam_loc522[14:0]) ? cam_loc522 : 11'd522 ) |
 ( (snoop_in == cam_loc523[14:0]) ? cam_loc523 : 11'd523 ) |
 ( (snoop_in == cam_loc524[14:0]) ? cam_loc524 : 11'd524 ) |
 ( (snoop_in == cam_loc525[14:0]) ? cam_loc525 : 11'd525 ) |
 ( (snoop_in == cam_loc526[14:0]) ? cam_loc526 : 11'd526 ) |
 ( (snoop_in == cam_loc527[14:0]) ? cam_loc527 : 11'd527 ) |
 ( (snoop_in == cam_loc528[14:0]) ? cam_loc528 : 11'd528 ) |
 ( (snoop_in == cam_loc529[14:0]) ? cam_loc529 : 11'd529 ) |
 ( (snoop_in == cam_loc530[14:0]) ? cam_loc530 : 11'd530 ) |
 ( (snoop_in == cam_loc531[14:0]) ? cam_loc531 : 11'd531 ) |
 ( (snoop_in == cam_loc532[14:0]) ? cam_loc532 : 11'd532 ) |
 ( (snoop_in == cam_loc533[14:0]) ? cam_loc533 : 11'd533 ) |
 ( (snoop_in == cam_loc534[14:0]) ? cam_loc534 : 11'd534 ) |
 ( (snoop_in == cam_loc535[14:0]) ? cam_loc535 : 11'd535 ) |
 ( (snoop_in == cam_loc536[14:0]) ? cam_loc536 : 11'd536 ) |
 ( (snoop_in == cam_loc537[14:0]) ? cam_loc537 : 11'd537 ) |
 ( (snoop_in == cam_loc538[14:0]) ? cam_loc538 : 11'd538 ) |
 ( (snoop_in == cam_loc539[14:0]) ? cam_loc539 : 11'd539 ) |
 ( (snoop_in == cam_loc540[14:0]) ? cam_loc540 : 11'd540 ) |
 ( (snoop_in == cam_loc541[14:0]) ? cam_loc541 : 11'd541 ) |
 ( (snoop_in == cam_loc542[14:0]) ? cam_loc542 : 11'd542 ) |
 ( (snoop_in == cam_loc543[14:0]) ? cam_loc543 : 11'd543 ) |
 ( (snoop_in == cam_loc544[14:0]) ? cam_loc544 : 11'd544 ) |
 ( (snoop_in == cam_loc545[14:0]) ? cam_loc545 : 11'd545 ) |
 ( (snoop_in == cam_loc546[14:0]) ? cam_loc546 : 11'd546 ) |
 ( (snoop_in == cam_loc547[14:0]) ? cam_loc547 : 11'd547 ) |
 ( (snoop_in == cam_loc548[14:0]) ? cam_loc548 : 11'd548 ) |
 ( (snoop_in == cam_loc549[14:0]) ? cam_loc549 : 11'd549 ) |
 ( (snoop_in == cam_loc550[14:0]) ? cam_loc550 : 11'd550 ) |
 ( (snoop_in == cam_loc551[14:0]) ? cam_loc551 : 11'd551 ) |
 ( (snoop_in == cam_loc552[14:0]) ? cam_loc552 : 11'd552 ) |
 ( (snoop_in == cam_loc553[14:0]) ? cam_loc553 : 11'd553 ) |
 ( (snoop_in == cam_loc554[14:0]) ? cam_loc554 : 11'd554 ) |
 ( (snoop_in == cam_loc555[14:0]) ? cam_loc555 : 11'd555 ) |
 ( (snoop_in == cam_loc556[14:0]) ? cam_loc556 : 11'd556 ) |
 ( (snoop_in == cam_loc557[14:0]) ? cam_loc557 : 11'd557 ) |
 ( (snoop_in == cam_loc558[14:0]) ? cam_loc558 : 11'd558 ) |
 ( (snoop_in == cam_loc559[14:0]) ? cam_loc559 : 11'd559 ) |
 ( (snoop_in == cam_loc560[14:0]) ? cam_loc560 : 11'd560 ) |
 ( (snoop_in == cam_loc561[14:0]) ? cam_loc561 : 11'd561 ) |
 ( (snoop_in == cam_loc562[14:0]) ? cam_loc562 : 11'd562 ) |
 ( (snoop_in == cam_loc563[14:0]) ? cam_loc563 : 11'd563 ) |
 ( (snoop_in == cam_loc564[14:0]) ? cam_loc564 : 11'd564 ) |
 ( (snoop_in == cam_loc565[14:0]) ? cam_loc565 : 11'd565 ) |
 ( (snoop_in == cam_loc566[14:0]) ? cam_loc566 : 11'd566 ) |
 ( (snoop_in == cam_loc567[14:0]) ? cam_loc567 : 11'd567 ) |
 ( (snoop_in == cam_loc568[14:0]) ? cam_loc568 : 11'd568 ) |
 ( (snoop_in == cam_loc569[14:0]) ? cam_loc569 : 11'd569 ) |
 ( (snoop_in == cam_loc570[14:0]) ? cam_loc570 : 11'd570 ) |
 ( (snoop_in == cam_loc571[14:0]) ? cam_loc571 : 11'd571 ) |
 ( (snoop_in == cam_loc572[14:0]) ? cam_loc572 : 11'd572 ) |
 ( (snoop_in == cam_loc573[14:0]) ? cam_loc573 : 11'd573 ) |
 ( (snoop_in == cam_loc574[14:0]) ? cam_loc574 : 11'd574 ) |
 ( (snoop_in == cam_loc575[14:0]) ? cam_loc575 : 11'd575 ) |
 ( (snoop_in == cam_loc576[14:0]) ? cam_loc576 : 11'd576 ) |
 ( (snoop_in == cam_loc577[14:0]) ? cam_loc577 : 11'd577 ) |
 ( (snoop_in == cam_loc578[14:0]) ? cam_loc578 : 11'd578 ) |
 ( (snoop_in == cam_loc579[14:0]) ? cam_loc579 : 11'd579 ) |
 ( (snoop_in == cam_loc580[14:0]) ? cam_loc580 : 11'd580 ) |
 ( (snoop_in == cam_loc581[14:0]) ? cam_loc581 : 11'd581 ) |
 ( (snoop_in == cam_loc582[14:0]) ? cam_loc582 : 11'd582 ) |
 ( (snoop_in == cam_loc583[14:0]) ? cam_loc583 : 11'd583 ) |
 ( (snoop_in == cam_loc584[14:0]) ? cam_loc584 : 11'd584 ) |
 ( (snoop_in == cam_loc585[14:0]) ? cam_loc585 : 11'd585 ) |
 ( (snoop_in == cam_loc586[14:0]) ? cam_loc586 : 11'd586 ) |
 ( (snoop_in == cam_loc587[14:0]) ? cam_loc587 : 11'd587 ) |
 ( (snoop_in == cam_loc588[14:0]) ? cam_loc588 : 11'd588 ) |
 ( (snoop_in == cam_loc589[14:0]) ? cam_loc589 : 11'd589 ) |
 ( (snoop_in == cam_loc590[14:0]) ? cam_loc590 : 11'd590 ) |
 ( (snoop_in == cam_loc591[14:0]) ? cam_loc591 : 11'd591 ) |
 ( (snoop_in == cam_loc592[14:0]) ? cam_loc592 : 11'd592 ) |
 ( (snoop_in == cam_loc593[14:0]) ? cam_loc593 : 11'd593 ) |
 ( (snoop_in == cam_loc594[14:0]) ? cam_loc594 : 11'd594 ) |
 ( (snoop_in == cam_loc595[14:0]) ? cam_loc595 : 11'd595 ) |
 ( (snoop_in == cam_loc596[14:0]) ? cam_loc596 : 11'd596 ) |
 ( (snoop_in == cam_loc597[14:0]) ? cam_loc597 : 11'd597 ) |
 ( (snoop_in == cam_loc598[14:0]) ? cam_loc598 : 11'd598 ) |
 ( (snoop_in == cam_loc599[14:0]) ? cam_loc599 : 11'd599 ) |
 ( (snoop_in == cam_loc600[14:0]) ? cam_loc600 : 11'd600 ) |
 ( (snoop_in == cam_loc601[14:0]) ? cam_loc601 : 11'd601 ) |
 ( (snoop_in == cam_loc602[14:0]) ? cam_loc602 : 11'd602 ) |
 ( (snoop_in == cam_loc603[14:0]) ? cam_loc603 : 11'd603 ) |
 ( (snoop_in == cam_loc604[14:0]) ? cam_loc604 : 11'd604 ) |
 ( (snoop_in == cam_loc605[14:0]) ? cam_loc605 : 11'd605 ) |
 ( (snoop_in == cam_loc606[14:0]) ? cam_loc606 : 11'd606 ) |
 ( (snoop_in == cam_loc607[14:0]) ? cam_loc607 : 11'd607 ) |
 ( (snoop_in == cam_loc608[14:0]) ? cam_loc608 : 11'd608 ) |
 ( (snoop_in == cam_loc609[14:0]) ? cam_loc609 : 11'd609 ) |
 ( (snoop_in == cam_loc610[14:0]) ? cam_loc610 : 11'd610 ) |
 ( (snoop_in == cam_loc611[14:0]) ? cam_loc611 : 11'd611 ) |
 ( (snoop_in == cam_loc612[14:0]) ? cam_loc612 : 11'd612 ) |
 ( (snoop_in == cam_loc613[14:0]) ? cam_loc613 : 11'd613 ) |
 ( (snoop_in == cam_loc614[14:0]) ? cam_loc614 : 11'd614 ) |
 ( (snoop_in == cam_loc615[14:0]) ? cam_loc615 : 11'd615 ) |
 ( (snoop_in == cam_loc616[14:0]) ? cam_loc616 : 11'd616 ) |
 ( (snoop_in == cam_loc617[14:0]) ? cam_loc617 : 11'd617 ) |
 ( (snoop_in == cam_loc618[14:0]) ? cam_loc618 : 11'd618 ) |
 ( (snoop_in == cam_loc619[14:0]) ? cam_loc619 : 11'd619 ) |
 ( (snoop_in == cam_loc620[14:0]) ? cam_loc620 : 11'd620 ) |
 ( (snoop_in == cam_loc621[14:0]) ? cam_loc621 : 11'd621 ) |
 ( (snoop_in == cam_loc622[14:0]) ? cam_loc622 : 11'd622 ) |
 ( (snoop_in == cam_loc623[14:0]) ? cam_loc623 : 11'd623 ) |
 ( (snoop_in == cam_loc624[14:0]) ? cam_loc624 : 11'd624 ) |
 ( (snoop_in == cam_loc625[14:0]) ? cam_loc625 : 11'd625 ) |
 ( (snoop_in == cam_loc626[14:0]) ? cam_loc626 : 11'd626 ) |
 ( (snoop_in == cam_loc627[14:0]) ? cam_loc627 : 11'd627 ) |
 ( (snoop_in == cam_loc628[14:0]) ? cam_loc628 : 11'd628 ) |
 ( (snoop_in == cam_loc629[14:0]) ? cam_loc629 : 11'd629 ) |
 ( (snoop_in == cam_loc630[14:0]) ? cam_loc630 : 11'd630 ) |
 ( (snoop_in == cam_loc631[14:0]) ? cam_loc631 : 11'd631 ) |
 ( (snoop_in == cam_loc632[14:0]) ? cam_loc632 : 11'd632 ) |
 ( (snoop_in == cam_loc633[14:0]) ? cam_loc633 : 11'd633 ) |
 ( (snoop_in == cam_loc634[14:0]) ? cam_loc634 : 11'd634 ) |
 ( (snoop_in == cam_loc635[14:0]) ? cam_loc635 : 11'd635 ) |
 ( (snoop_in == cam_loc636[14:0]) ? cam_loc636 : 11'd636 ) |
 ( (snoop_in == cam_loc637[14:0]) ? cam_loc637 : 11'd637 ) |
 ( (snoop_in == cam_loc638[14:0]) ? cam_loc638 : 11'd638 ) |
 ( (snoop_in == cam_loc639[14:0]) ? cam_loc639 : 11'd639 ) |
 ( (snoop_in == cam_loc640[14:0]) ? cam_loc640 : 11'd640 ) |
 ( (snoop_in == cam_loc641[14:0]) ? cam_loc641 : 11'd641 ) |
 ( (snoop_in == cam_loc642[14:0]) ? cam_loc642 : 11'd642 ) |
 ( (snoop_in == cam_loc643[14:0]) ? cam_loc643 : 11'd643 ) |
 ( (snoop_in == cam_loc644[14:0]) ? cam_loc644 : 11'd644 ) |
 ( (snoop_in == cam_loc645[14:0]) ? cam_loc645 : 11'd645 ) |
 ( (snoop_in == cam_loc646[14:0]) ? cam_loc646 : 11'd646 ) |
 ( (snoop_in == cam_loc647[14:0]) ? cam_loc647 : 11'd647 ) |
 ( (snoop_in == cam_loc648[14:0]) ? cam_loc648 : 11'd648 ) |
 ( (snoop_in == cam_loc649[14:0]) ? cam_loc649 : 11'd649 ) |
 ( (snoop_in == cam_loc650[14:0]) ? cam_loc650 : 11'd650 ) |
 ( (snoop_in == cam_loc651[14:0]) ? cam_loc651 : 11'd651 ) |
 ( (snoop_in == cam_loc652[14:0]) ? cam_loc652 : 11'd652 ) |
 ( (snoop_in == cam_loc653[14:0]) ? cam_loc653 : 11'd653 ) |
 ( (snoop_in == cam_loc654[14:0]) ? cam_loc654 : 11'd654 ) |
 ( (snoop_in == cam_loc655[14:0]) ? cam_loc655 : 11'd655 ) |
 ( (snoop_in == cam_loc656[14:0]) ? cam_loc656 : 11'd656 ) |
 ( (snoop_in == cam_loc657[14:0]) ? cam_loc657 : 11'd657 ) |
 ( (snoop_in == cam_loc658[14:0]) ? cam_loc658 : 11'd658 ) |
 ( (snoop_in == cam_loc659[14:0]) ? cam_loc659 : 11'd659 ) |
 ( (snoop_in == cam_loc660[14:0]) ? cam_loc660 : 11'd660 ) |
 ( (snoop_in == cam_loc661[14:0]) ? cam_loc661 : 11'd661 ) |
 ( (snoop_in == cam_loc662[14:0]) ? cam_loc662 : 11'd662 ) |
 ( (snoop_in == cam_loc663[14:0]) ? cam_loc663 : 11'd663 ) |
 ( (snoop_in == cam_loc664[14:0]) ? cam_loc664 : 11'd664 ) |
 ( (snoop_in == cam_loc665[14:0]) ? cam_loc665 : 11'd665 ) |
 ( (snoop_in == cam_loc666[14:0]) ? cam_loc666 : 11'd666 ) |
 ( (snoop_in == cam_loc667[14:0]) ? cam_loc667 : 11'd667 ) |
 ( (snoop_in == cam_loc668[14:0]) ? cam_loc668 : 11'd668 ) |
 ( (snoop_in == cam_loc669[14:0]) ? cam_loc669 : 11'd669 ) |
 ( (snoop_in == cam_loc670[14:0]) ? cam_loc670 : 11'd670 ) |
 ( (snoop_in == cam_loc671[14:0]) ? cam_loc671 : 11'd671 ) |
 ( (snoop_in == cam_loc672[14:0]) ? cam_loc672 : 11'd672 ) |
 ( (snoop_in == cam_loc673[14:0]) ? cam_loc673 : 11'd673 ) |
 ( (snoop_in == cam_loc674[14:0]) ? cam_loc674 : 11'd674 ) |
 ( (snoop_in == cam_loc675[14:0]) ? cam_loc675 : 11'd675 ) |
 ( (snoop_in == cam_loc676[14:0]) ? cam_loc676 : 11'd676 ) |
 ( (snoop_in == cam_loc677[14:0]) ? cam_loc677 : 11'd677 ) |
 ( (snoop_in == cam_loc678[14:0]) ? cam_loc678 : 11'd678 ) |
 ( (snoop_in == cam_loc679[14:0]) ? cam_loc679 : 11'd679 ) |
 ( (snoop_in == cam_loc680[14:0]) ? cam_loc680 : 11'd680 ) |
 ( (snoop_in == cam_loc681[14:0]) ? cam_loc681 : 11'd681 ) |
 ( (snoop_in == cam_loc682[14:0]) ? cam_loc682 : 11'd682 ) |
 ( (snoop_in == cam_loc683[14:0]) ? cam_loc683 : 11'd683 ) |
 ( (snoop_in == cam_loc684[14:0]) ? cam_loc684 : 11'd684 ) |
 ( (snoop_in == cam_loc685[14:0]) ? cam_loc685 : 11'd685 ) |
 ( (snoop_in == cam_loc686[14:0]) ? cam_loc686 : 11'd686 ) |
 ( (snoop_in == cam_loc687[14:0]) ? cam_loc687 : 11'd687 ) |
 ( (snoop_in == cam_loc688[14:0]) ? cam_loc688 : 11'd688 ) |
 ( (snoop_in == cam_loc689[14:0]) ? cam_loc689 : 11'd689 ) |
 ( (snoop_in == cam_loc690[14:0]) ? cam_loc690 : 11'd690 ) |
 ( (snoop_in == cam_loc691[14:0]) ? cam_loc691 : 11'd691 ) |
 ( (snoop_in == cam_loc692[14:0]) ? cam_loc692 : 11'd692 ) |
 ( (snoop_in == cam_loc693[14:0]) ? cam_loc693 : 11'd693 ) |
 ( (snoop_in == cam_loc694[14:0]) ? cam_loc694 : 11'd694 ) |
 ( (snoop_in == cam_loc695[14:0]) ? cam_loc695 : 11'd695 ) |
 ( (snoop_in == cam_loc696[14:0]) ? cam_loc696 : 11'd696 ) |
 ( (snoop_in == cam_loc697[14:0]) ? cam_loc697 : 11'd697 ) |
 ( (snoop_in == cam_loc698[14:0]) ? cam_loc698 : 11'd698 ) |
 ( (snoop_in == cam_loc699[14:0]) ? cam_loc699 : 11'd699 ) |
 ( (snoop_in == cam_loc700[14:0]) ? cam_loc700 : 11'd700 ) |
 ( (snoop_in == cam_loc701[14:0]) ? cam_loc701 : 11'd701 ) |
 ( (snoop_in == cam_loc702[14:0]) ? cam_loc702 : 11'd702 ) |
 ( (snoop_in == cam_loc703[14:0]) ? cam_loc703 : 11'd703 ) |
 ( (snoop_in == cam_loc704[14:0]) ? cam_loc704 : 11'd704 ) |
 ( (snoop_in == cam_loc705[14:0]) ? cam_loc705 : 11'd705 ) |
 ( (snoop_in == cam_loc706[14:0]) ? cam_loc706 : 11'd706 ) |
 ( (snoop_in == cam_loc707[14:0]) ? cam_loc707 : 11'd707 ) |
 ( (snoop_in == cam_loc708[14:0]) ? cam_loc708 : 11'd708 ) |
 ( (snoop_in == cam_loc709[14:0]) ? cam_loc709 : 11'd709 ) |
 ( (snoop_in == cam_loc710[14:0]) ? cam_loc710 : 11'd710 ) |
 ( (snoop_in == cam_loc711[14:0]) ? cam_loc711 : 11'd711 ) |
 ( (snoop_in == cam_loc712[14:0]) ? cam_loc712 : 11'd712 ) |
 ( (snoop_in == cam_loc713[14:0]) ? cam_loc713 : 11'd713 ) |
 ( (snoop_in == cam_loc714[14:0]) ? cam_loc714 : 11'd714 ) |
 ( (snoop_in == cam_loc715[14:0]) ? cam_loc715 : 11'd715 ) |
 ( (snoop_in == cam_loc716[14:0]) ? cam_loc716 : 11'd716 ) |
 ( (snoop_in == cam_loc717[14:0]) ? cam_loc717 : 11'd717 ) |
 ( (snoop_in == cam_loc718[14:0]) ? cam_loc718 : 11'd718 ) |
 ( (snoop_in == cam_loc719[14:0]) ? cam_loc719 : 11'd719 ) |
 ( (snoop_in == cam_loc720[14:0]) ? cam_loc720 : 11'd720 ) |
 ( (snoop_in == cam_loc721[14:0]) ? cam_loc721 : 11'd721 ) |
 ( (snoop_in == cam_loc722[14:0]) ? cam_loc722 : 11'd722 ) |
 ( (snoop_in == cam_loc723[14:0]) ? cam_loc723 : 11'd723 ) |
 ( (snoop_in == cam_loc724[14:0]) ? cam_loc724 : 11'd724 ) |
 ( (snoop_in == cam_loc725[14:0]) ? cam_loc725 : 11'd725 ) |
 ( (snoop_in == cam_loc726[14:0]) ? cam_loc726 : 11'd726 ) |
 ( (snoop_in == cam_loc727[14:0]) ? cam_loc727 : 11'd727 ) |
 ( (snoop_in == cam_loc728[14:0]) ? cam_loc728 : 11'd728 ) |
 ( (snoop_in == cam_loc729[14:0]) ? cam_loc729 : 11'd729 ) |
 ( (snoop_in == cam_loc730[14:0]) ? cam_loc730 : 11'd730 ) |
 ( (snoop_in == cam_loc731[14:0]) ? cam_loc731 : 11'd731 ) |
 ( (snoop_in == cam_loc732[14:0]) ? cam_loc732 : 11'd732 ) |
 ( (snoop_in == cam_loc733[14:0]) ? cam_loc733 : 11'd733 ) |
 ( (snoop_in == cam_loc734[14:0]) ? cam_loc734 : 11'd734 ) |
 ( (snoop_in == cam_loc735[14:0]) ? cam_loc735 : 11'd735 ) |
 ( (snoop_in == cam_loc736[14:0]) ? cam_loc736 : 11'd736 ) |
 ( (snoop_in == cam_loc737[14:0]) ? cam_loc737 : 11'd737 ) |
 ( (snoop_in == cam_loc738[14:0]) ? cam_loc738 : 11'd738 ) |
 ( (snoop_in == cam_loc739[14:0]) ? cam_loc739 : 11'd739 ) |
 ( (snoop_in == cam_loc740[14:0]) ? cam_loc740 : 11'd740 ) |
 ( (snoop_in == cam_loc741[14:0]) ? cam_loc741 : 11'd741 ) |
 ( (snoop_in == cam_loc742[14:0]) ? cam_loc742 : 11'd742 ) |
 ( (snoop_in == cam_loc743[14:0]) ? cam_loc743 : 11'd743 ) |
 ( (snoop_in == cam_loc744[14:0]) ? cam_loc744 : 11'd744 ) |
 ( (snoop_in == cam_loc745[14:0]) ? cam_loc745 : 11'd745 ) |
 ( (snoop_in == cam_loc746[14:0]) ? cam_loc746 : 11'd746 ) |
 ( (snoop_in == cam_loc747[14:0]) ? cam_loc747 : 11'd747 ) |
 ( (snoop_in == cam_loc748[14:0]) ? cam_loc748 : 11'd748 ) |
 ( (snoop_in == cam_loc749[14:0]) ? cam_loc749 : 11'd749 ) |
 ( (snoop_in == cam_loc750[14:0]) ? cam_loc750 : 11'd750 ) |
 ( (snoop_in == cam_loc751[14:0]) ? cam_loc751 : 11'd751 ) |
 ( (snoop_in == cam_loc752[14:0]) ? cam_loc752 : 11'd752 ) |
 ( (snoop_in == cam_loc753[14:0]) ? cam_loc753 : 11'd753 ) |
 ( (snoop_in == cam_loc754[14:0]) ? cam_loc754 : 11'd754 ) |
 ( (snoop_in == cam_loc755[14:0]) ? cam_loc755 : 11'd755 ) |
 ( (snoop_in == cam_loc756[14:0]) ? cam_loc756 : 11'd756 ) |
 ( (snoop_in == cam_loc757[14:0]) ? cam_loc757 : 11'd757 ) |
 ( (snoop_in == cam_loc758[14:0]) ? cam_loc758 : 11'd758 ) |
 ( (snoop_in == cam_loc759[14:0]) ? cam_loc759 : 11'd759 ) |
 ( (snoop_in == cam_loc760[14:0]) ? cam_loc760 : 11'd760 ) |
 ( (snoop_in == cam_loc761[14:0]) ? cam_loc761 : 11'd761 ) |
 ( (snoop_in == cam_loc762[14:0]) ? cam_loc762 : 11'd762 ) |
 ( (snoop_in == cam_loc763[14:0]) ? cam_loc763 : 11'd763 ) |
 ( (snoop_in == cam_loc764[14:0]) ? cam_loc764 : 11'd764 ) |
 ( (snoop_in == cam_loc765[14:0]) ? cam_loc765 : 11'd765 ) |
 ( (snoop_in == cam_loc766[14:0]) ? cam_loc766 : 11'd766 ) |
 ( (snoop_in == cam_loc767[14:0]) ? cam_loc767 : 11'd767 ) |
 ( (snoop_in == cam_loc768[14:0]) ? cam_loc768 : 11'd768 ) |
 ( (snoop_in == cam_loc769[14:0]) ? cam_loc769 : 11'd769 ) |
 ( (snoop_in == cam_loc770[14:0]) ? cam_loc770 : 11'd770 ) |
 ( (snoop_in == cam_loc771[14:0]) ? cam_loc771 : 11'd771 ) |
 ( (snoop_in == cam_loc772[14:0]) ? cam_loc772 : 11'd772 ) |
 ( (snoop_in == cam_loc773[14:0]) ? cam_loc773 : 11'd773 ) |
 ( (snoop_in == cam_loc774[14:0]) ? cam_loc774 : 11'd774 ) |
 ( (snoop_in == cam_loc775[14:0]) ? cam_loc775 : 11'd775 ) |
 ( (snoop_in == cam_loc776[14:0]) ? cam_loc776 : 11'd776 ) |
 ( (snoop_in == cam_loc777[14:0]) ? cam_loc777 : 11'd777 ) |
 ( (snoop_in == cam_loc778[14:0]) ? cam_loc778 : 11'd778 ) |
 ( (snoop_in == cam_loc779[14:0]) ? cam_loc779 : 11'd779 ) |
 ( (snoop_in == cam_loc780[14:0]) ? cam_loc780 : 11'd780 ) |
 ( (snoop_in == cam_loc781[14:0]) ? cam_loc781 : 11'd781 ) |
 ( (snoop_in == cam_loc782[14:0]) ? cam_loc782 : 11'd782 ) |
 ( (snoop_in == cam_loc783[14:0]) ? cam_loc783 : 11'd783 ) |
 ( (snoop_in == cam_loc784[14:0]) ? cam_loc784 : 11'd784 ) |
 ( (snoop_in == cam_loc785[14:0]) ? cam_loc785 : 11'd785 ) |
 ( (snoop_in == cam_loc786[14:0]) ? cam_loc786 : 11'd786 ) |
 ( (snoop_in == cam_loc787[14:0]) ? cam_loc787 : 11'd787 ) |
 ( (snoop_in == cam_loc788[14:0]) ? cam_loc788 : 11'd788 ) |
 ( (snoop_in == cam_loc789[14:0]) ? cam_loc789 : 11'd789 ) |
 ( (snoop_in == cam_loc790[14:0]) ? cam_loc790 : 11'd790 ) |
 ( (snoop_in == cam_loc791[14:0]) ? cam_loc791 : 11'd791 ) |
 ( (snoop_in == cam_loc792[14:0]) ? cam_loc792 : 11'd792 ) |
 ( (snoop_in == cam_loc793[14:0]) ? cam_loc793 : 11'd793 ) |
 ( (snoop_in == cam_loc794[14:0]) ? cam_loc794 : 11'd794 ) |
 ( (snoop_in == cam_loc795[14:0]) ? cam_loc795 : 11'd795 ) |
 ( (snoop_in == cam_loc796[14:0]) ? cam_loc796 : 11'd796 ) |
 ( (snoop_in == cam_loc797[14:0]) ? cam_loc797 : 11'd797 ) |
 ( (snoop_in == cam_loc798[14:0]) ? cam_loc798 : 11'd798 ) |
 ( (snoop_in == cam_loc799[14:0]) ? cam_loc799 : 11'd799 ) |
 ( (snoop_in == cam_loc800[14:0]) ? cam_loc800 : 11'd800 ) |
 ( (snoop_in == cam_loc801[14:0]) ? cam_loc801 : 11'd801 ) |
 ( (snoop_in == cam_loc802[14:0]) ? cam_loc802 : 11'd802 ) |
 ( (snoop_in == cam_loc803[14:0]) ? cam_loc803 : 11'd803 ) |
 ( (snoop_in == cam_loc804[14:0]) ? cam_loc804 : 11'd804 ) |
 ( (snoop_in == cam_loc805[14:0]) ? cam_loc805 : 11'd805 ) |
 ( (snoop_in == cam_loc806[14:0]) ? cam_loc806 : 11'd806 ) |
 ( (snoop_in == cam_loc807[14:0]) ? cam_loc807 : 11'd807 ) |
 ( (snoop_in == cam_loc808[14:0]) ? cam_loc808 : 11'd808 ) |
 ( (snoop_in == cam_loc809[14:0]) ? cam_loc809 : 11'd809 ) |
 ( (snoop_in == cam_loc810[14:0]) ? cam_loc810 : 11'd810 ) |
 ( (snoop_in == cam_loc811[14:0]) ? cam_loc811 : 11'd811 ) |
 ( (snoop_in == cam_loc812[14:0]) ? cam_loc812 : 11'd812 ) |
 ( (snoop_in == cam_loc813[14:0]) ? cam_loc813 : 11'd813 ) |
 ( (snoop_in == cam_loc814[14:0]) ? cam_loc814 : 11'd814 ) |
 ( (snoop_in == cam_loc815[14:0]) ? cam_loc815 : 11'd815 ) |
 ( (snoop_in == cam_loc816[14:0]) ? cam_loc816 : 11'd816 ) |
 ( (snoop_in == cam_loc817[14:0]) ? cam_loc817 : 11'd817 ) |
 ( (snoop_in == cam_loc818[14:0]) ? cam_loc818 : 11'd818 ) |
 ( (snoop_in == cam_loc819[14:0]) ? cam_loc819 : 11'd819 ) |
 ( (snoop_in == cam_loc820[14:0]) ? cam_loc820 : 11'd820 ) |
 ( (snoop_in == cam_loc821[14:0]) ? cam_loc821 : 11'd821 ) |
 ( (snoop_in == cam_loc822[14:0]) ? cam_loc822 : 11'd822 ) |
 ( (snoop_in == cam_loc823[14:0]) ? cam_loc823 : 11'd823 ) |
 ( (snoop_in == cam_loc824[14:0]) ? cam_loc824 : 11'd824 ) |
 ( (snoop_in == cam_loc825[14:0]) ? cam_loc825 : 11'd825 ) |
 ( (snoop_in == cam_loc826[14:0]) ? cam_loc826 : 11'd826 ) |
 ( (snoop_in == cam_loc827[14:0]) ? cam_loc827 : 11'd827 ) |
 ( (snoop_in == cam_loc828[14:0]) ? cam_loc828 : 11'd828 ) |
 ( (snoop_in == cam_loc829[14:0]) ? cam_loc829 : 11'd829 ) |
 ( (snoop_in == cam_loc830[14:0]) ? cam_loc830 : 11'd830 ) |
 ( (snoop_in == cam_loc831[14:0]) ? cam_loc831 : 11'd831 ) |
 ( (snoop_in == cam_loc832[14:0]) ? cam_loc832 : 11'd832 ) |
 ( (snoop_in == cam_loc833[14:0]) ? cam_loc833 : 11'd833 ) |
 ( (snoop_in == cam_loc834[14:0]) ? cam_loc834 : 11'd834 ) |
 ( (snoop_in == cam_loc835[14:0]) ? cam_loc835 : 11'd835 ) |
 ( (snoop_in == cam_loc836[14:0]) ? cam_loc836 : 11'd836 ) |
 ( (snoop_in == cam_loc837[14:0]) ? cam_loc837 : 11'd837 ) |
 ( (snoop_in == cam_loc838[14:0]) ? cam_loc838 : 11'd838 ) |
 ( (snoop_in == cam_loc839[14:0]) ? cam_loc839 : 11'd839 ) |
 ( (snoop_in == cam_loc840[14:0]) ? cam_loc840 : 11'd840 ) |
 ( (snoop_in == cam_loc841[14:0]) ? cam_loc841 : 11'd841 ) |
 ( (snoop_in == cam_loc842[14:0]) ? cam_loc842 : 11'd842 ) |
 ( (snoop_in == cam_loc843[14:0]) ? cam_loc843 : 11'd843 ) |
 ( (snoop_in == cam_loc844[14:0]) ? cam_loc844 : 11'd844 ) |
 ( (snoop_in == cam_loc845[14:0]) ? cam_loc845 : 11'd845 ) |
 ( (snoop_in == cam_loc846[14:0]) ? cam_loc846 : 11'd846 ) |
 ( (snoop_in == cam_loc847[14:0]) ? cam_loc847 : 11'd847 ) |
 ( (snoop_in == cam_loc848[14:0]) ? cam_loc848 : 11'd848 ) |
 ( (snoop_in == cam_loc849[14:0]) ? cam_loc849 : 11'd849 ) |
 ( (snoop_in == cam_loc850[14:0]) ? cam_loc850 : 11'd850 ) |
 ( (snoop_in == cam_loc851[14:0]) ? cam_loc851 : 11'd851 ) |
 ( (snoop_in == cam_loc852[14:0]) ? cam_loc852 : 11'd852 ) |
 ( (snoop_in == cam_loc853[14:0]) ? cam_loc853 : 11'd853 ) |
 ( (snoop_in == cam_loc854[14:0]) ? cam_loc854 : 11'd854 ) |
 ( (snoop_in == cam_loc855[14:0]) ? cam_loc855 : 11'd855 ) |
 ( (snoop_in == cam_loc856[14:0]) ? cam_loc856 : 11'd856 ) |
 ( (snoop_in == cam_loc857[14:0]) ? cam_loc857 : 11'd857 ) |
 ( (snoop_in == cam_loc858[14:0]) ? cam_loc858 : 11'd858 ) |
 ( (snoop_in == cam_loc859[14:0]) ? cam_loc859 : 11'd859 ) |
 ( (snoop_in == cam_loc860[14:0]) ? cam_loc860 : 11'd860 ) |
 ( (snoop_in == cam_loc861[14:0]) ? cam_loc861 : 11'd861 ) |
 ( (snoop_in == cam_loc862[14:0]) ? cam_loc862 : 11'd862 ) |
 ( (snoop_in == cam_loc863[14:0]) ? cam_loc863 : 11'd863 ) |
 ( (snoop_in == cam_loc864[14:0]) ? cam_loc864 : 11'd864 ) |
 ( (snoop_in == cam_loc865[14:0]) ? cam_loc865 : 11'd865 ) |
 ( (snoop_in == cam_loc866[14:0]) ? cam_loc866 : 11'd866 ) |
 ( (snoop_in == cam_loc867[14:0]) ? cam_loc867 : 11'd867 ) |
 ( (snoop_in == cam_loc868[14:0]) ? cam_loc868 : 11'd868 ) |
 ( (snoop_in == cam_loc869[14:0]) ? cam_loc869 : 11'd869 ) |
 ( (snoop_in == cam_loc870[14:0]) ? cam_loc870 : 11'd870 ) |
 ( (snoop_in == cam_loc871[14:0]) ? cam_loc871 : 11'd871 ) |
 ( (snoop_in == cam_loc872[14:0]) ? cam_loc872 : 11'd872 ) |
 ( (snoop_in == cam_loc873[14:0]) ? cam_loc873 : 11'd873 ) |
 ( (snoop_in == cam_loc874[14:0]) ? cam_loc874 : 11'd874 ) |
 ( (snoop_in == cam_loc875[14:0]) ? cam_loc875 : 11'd875 ) |
 ( (snoop_in == cam_loc876[14:0]) ? cam_loc876 : 11'd876 ) |
 ( (snoop_in == cam_loc877[14:0]) ? cam_loc877 : 11'd877 ) |
 ( (snoop_in == cam_loc878[14:0]) ? cam_loc878 : 11'd878 ) |
 ( (snoop_in == cam_loc879[14:0]) ? cam_loc879 : 11'd879 ) |
 ( (snoop_in == cam_loc880[14:0]) ? cam_loc880 : 11'd880 ) |
 ( (snoop_in == cam_loc881[14:0]) ? cam_loc881 : 11'd881 ) |
 ( (snoop_in == cam_loc882[14:0]) ? cam_loc882 : 11'd882 ) |
 ( (snoop_in == cam_loc883[14:0]) ? cam_loc883 : 11'd883 ) |
 ( (snoop_in == cam_loc884[14:0]) ? cam_loc884 : 11'd884 ) |
 ( (snoop_in == cam_loc885[14:0]) ? cam_loc885 : 11'd885 ) |
 ( (snoop_in == cam_loc886[14:0]) ? cam_loc886 : 11'd886 ) |
 ( (snoop_in == cam_loc887[14:0]) ? cam_loc887 : 11'd887 ) |
 ( (snoop_in == cam_loc888[14:0]) ? cam_loc888 : 11'd888 ) |
 ( (snoop_in == cam_loc889[14:0]) ? cam_loc889 : 11'd889 ) |
 ( (snoop_in == cam_loc890[14:0]) ? cam_loc890 : 11'd890 ) |
 ( (snoop_in == cam_loc891[14:0]) ? cam_loc891 : 11'd891 ) |
 ( (snoop_in == cam_loc892[14:0]) ? cam_loc892 : 11'd892 ) |
 ( (snoop_in == cam_loc893[14:0]) ? cam_loc893 : 11'd893 ) |
 ( (snoop_in == cam_loc894[14:0]) ? cam_loc894 : 11'd894 ) |
 ( (snoop_in == cam_loc895[14:0]) ? cam_loc895 : 11'd895 ) |
 ( (snoop_in == cam_loc896[14:0]) ? cam_loc896 : 11'd896 ) |
 ( (snoop_in == cam_loc897[14:0]) ? cam_loc897 : 11'd897 ) |
 ( (snoop_in == cam_loc898[14:0]) ? cam_loc898 : 11'd898 ) |
 ( (snoop_in == cam_loc899[14:0]) ? cam_loc899 : 11'd899 ) |
 ( (snoop_in == cam_loc900[14:0]) ? cam_loc900 : 11'd900 ) |
 ( (snoop_in == cam_loc901[14:0]) ? cam_loc901 : 11'd901 ) |
 ( (snoop_in == cam_loc902[14:0]) ? cam_loc902 : 11'd902 ) |
 ( (snoop_in == cam_loc903[14:0]) ? cam_loc903 : 11'd903 ) |
 ( (snoop_in == cam_loc904[14:0]) ? cam_loc904 : 11'd904 ) |
 ( (snoop_in == cam_loc905[14:0]) ? cam_loc905 : 11'd905 ) |
 ( (snoop_in == cam_loc906[14:0]) ? cam_loc906 : 11'd906 ) |
 ( (snoop_in == cam_loc907[14:0]) ? cam_loc907 : 11'd907 ) |
 ( (snoop_in == cam_loc908[14:0]) ? cam_loc908 : 11'd908 ) |
 ( (snoop_in == cam_loc909[14:0]) ? cam_loc909 : 11'd909 ) |
 ( (snoop_in == cam_loc910[14:0]) ? cam_loc910 : 11'd910 ) |
 ( (snoop_in == cam_loc911[14:0]) ? cam_loc911 : 11'd911 ) |
 ( (snoop_in == cam_loc912[14:0]) ? cam_loc912 : 11'd912 ) |
 ( (snoop_in == cam_loc913[14:0]) ? cam_loc913 : 11'd913 ) |
 ( (snoop_in == cam_loc914[14:0]) ? cam_loc914 : 11'd914 ) |
 ( (snoop_in == cam_loc915[14:0]) ? cam_loc915 : 11'd915 ) |
 ( (snoop_in == cam_loc916[14:0]) ? cam_loc916 : 11'd916 ) |
 ( (snoop_in == cam_loc917[14:0]) ? cam_loc917 : 11'd917 ) |
 ( (snoop_in == cam_loc918[14:0]) ? cam_loc918 : 11'd918 ) |
 ( (snoop_in == cam_loc919[14:0]) ? cam_loc919 : 11'd919 ) |
 ( (snoop_in == cam_loc920[14:0]) ? cam_loc920 : 11'd920 ) |
 ( (snoop_in == cam_loc921[14:0]) ? cam_loc921 : 11'd921 ) |
 ( (snoop_in == cam_loc922[14:0]) ? cam_loc922 : 11'd922 ) |
 ( (snoop_in == cam_loc923[14:0]) ? cam_loc923 : 11'd923 ) |
 ( (snoop_in == cam_loc924[14:0]) ? cam_loc924 : 11'd924 ) |
 ( (snoop_in == cam_loc925[14:0]) ? cam_loc925 : 11'd925 ) |
 ( (snoop_in == cam_loc926[14:0]) ? cam_loc926 : 11'd926 ) |
 ( (snoop_in == cam_loc927[14:0]) ? cam_loc927 : 11'd927 ) |
 ( (snoop_in == cam_loc928[14:0]) ? cam_loc928 : 11'd928 ) |
 ( (snoop_in == cam_loc929[14:0]) ? cam_loc929 : 11'd929 ) |
 ( (snoop_in == cam_loc930[14:0]) ? cam_loc930 : 11'd930 ) |
 ( (snoop_in == cam_loc931[14:0]) ? cam_loc931 : 11'd931 ) |
 ( (snoop_in == cam_loc932[14:0]) ? cam_loc932 : 11'd932 ) |
 ( (snoop_in == cam_loc933[14:0]) ? cam_loc933 : 11'd933 ) |
 ( (snoop_in == cam_loc934[14:0]) ? cam_loc934 : 11'd934 ) |
 ( (snoop_in == cam_loc935[14:0]) ? cam_loc935 : 11'd935 ) |
 ( (snoop_in == cam_loc936[14:0]) ? cam_loc936 : 11'd936 ) |
 ( (snoop_in == cam_loc937[14:0]) ? cam_loc937 : 11'd937 ) |
 ( (snoop_in == cam_loc938[14:0]) ? cam_loc938 : 11'd938 ) |
 ( (snoop_in == cam_loc939[14:0]) ? cam_loc939 : 11'd939 ) |
 ( (snoop_in == cam_loc940[14:0]) ? cam_loc940 : 11'd940 ) |
 ( (snoop_in == cam_loc941[14:0]) ? cam_loc941 : 11'd941 ) |
 ( (snoop_in == cam_loc942[14:0]) ? cam_loc942 : 11'd942 ) |
 ( (snoop_in == cam_loc943[14:0]) ? cam_loc943 : 11'd943 ) |
 ( (snoop_in == cam_loc944[14:0]) ? cam_loc944 : 11'd944 ) |
 ( (snoop_in == cam_loc945[14:0]) ? cam_loc945 : 11'd945 ) |
 ( (snoop_in == cam_loc946[14:0]) ? cam_loc946 : 11'd946 ) |
 ( (snoop_in == cam_loc947[14:0]) ? cam_loc947 : 11'd947 ) |
 ( (snoop_in == cam_loc948[14:0]) ? cam_loc948 : 11'd948 ) |
 ( (snoop_in == cam_loc949[14:0]) ? cam_loc949 : 11'd949 ) |
 ( (snoop_in == cam_loc950[14:0]) ? cam_loc950 : 11'd950 ) |
 ( (snoop_in == cam_loc951[14:0]) ? cam_loc951 : 11'd951 ) |
 ( (snoop_in == cam_loc952[14:0]) ? cam_loc952 : 11'd952 ) |
 ( (snoop_in == cam_loc953[14:0]) ? cam_loc953 : 11'd953 ) |
 ( (snoop_in == cam_loc954[14:0]) ? cam_loc954 : 11'd954 ) |
 ( (snoop_in == cam_loc955[14:0]) ? cam_loc955 : 11'd955 ) |
 ( (snoop_in == cam_loc956[14:0]) ? cam_loc956 : 11'd956 ) |
 ( (snoop_in == cam_loc957[14:0]) ? cam_loc957 : 11'd957 ) |
 ( (snoop_in == cam_loc958[14:0]) ? cam_loc958 : 11'd958 ) |
 ( (snoop_in == cam_loc959[14:0]) ? cam_loc959 : 11'd959 ) |
 ( (snoop_in == cam_loc960[14:0]) ? cam_loc960 : 11'd960 ) |
 ( (snoop_in == cam_loc961[14:0]) ? cam_loc961 : 11'd961 ) |
 ( (snoop_in == cam_loc962[14:0]) ? cam_loc962 : 11'd962 ) |
 ( (snoop_in == cam_loc963[14:0]) ? cam_loc963 : 11'd963 ) |
 ( (snoop_in == cam_loc964[14:0]) ? cam_loc964 : 11'd964 ) |
 ( (snoop_in == cam_loc965[14:0]) ? cam_loc965 : 11'd965 ) |
 ( (snoop_in == cam_loc966[14:0]) ? cam_loc966 : 11'd966 ) |
 ( (snoop_in == cam_loc967[14:0]) ? cam_loc967 : 11'd967 ) |
 ( (snoop_in == cam_loc968[14:0]) ? cam_loc968 : 11'd968 ) |
 ( (snoop_in == cam_loc969[14:0]) ? cam_loc969 : 11'd969 ) |
 ( (snoop_in == cam_loc970[14:0]) ? cam_loc970 : 11'd970 ) |
 ( (snoop_in == cam_loc971[14:0]) ? cam_loc971 : 11'd971 ) |
 ( (snoop_in == cam_loc972[14:0]) ? cam_loc972 : 11'd972 ) |
 ( (snoop_in == cam_loc973[14:0]) ? cam_loc973 : 11'd973 ) |
 ( (snoop_in == cam_loc974[14:0]) ? cam_loc974 : 11'd974 ) |
 ( (snoop_in == cam_loc975[14:0]) ? cam_loc975 : 11'd975 ) |
 ( (snoop_in == cam_loc976[14:0]) ? cam_loc976 : 11'd976 ) |
 ( (snoop_in == cam_loc977[14:0]) ? cam_loc977 : 11'd977 ) |
 ( (snoop_in == cam_loc978[14:0]) ? cam_loc978 : 11'd978 ) |
 ( (snoop_in == cam_loc979[14:0]) ? cam_loc979 : 11'd979 ) |
 ( (snoop_in == cam_loc980[14:0]) ? cam_loc980 : 11'd980 ) |
 ( (snoop_in == cam_loc981[14:0]) ? cam_loc981 : 11'd981 ) |
 ( (snoop_in == cam_loc982[14:0]) ? cam_loc982 : 11'd982 ) |
 ( (snoop_in == cam_loc983[14:0]) ? cam_loc983 : 11'd983 ) |
 ( (snoop_in == cam_loc984[14:0]) ? cam_loc984 : 11'd984 ) |
 ( (snoop_in == cam_loc985[14:0]) ? cam_loc985 : 11'd985 ) |
 ( (snoop_in == cam_loc986[14:0]) ? cam_loc986 : 11'd986 ) |
 ( (snoop_in == cam_loc987[14:0]) ? cam_loc987 : 11'd987 ) |
 ( (snoop_in == cam_loc988[14:0]) ? cam_loc988 : 11'd988 ) |
 ( (snoop_in == cam_loc989[14:0]) ? cam_loc989 : 11'd989 ) |
 ( (snoop_in == cam_loc990[14:0]) ? cam_loc990 : 11'd990 ) |
 ( (snoop_in == cam_loc991[14:0]) ? cam_loc991 : 11'd991 ) |
 ( (snoop_in == cam_loc992[14:0]) ? cam_loc992 : 11'd992 ) |
 ( (snoop_in == cam_loc993[14:0]) ? cam_loc993 : 11'd993 ) |
 ( (snoop_in == cam_loc994[14:0]) ? cam_loc994 : 11'd994 ) |
 ( (snoop_in == cam_loc995[14:0]) ? cam_loc995 : 11'd995 ) |
 ( (snoop_in == cam_loc996[14:0]) ? cam_loc996 : 11'd996 ) |
 ( (snoop_in == cam_loc997[14:0]) ? cam_loc997 : 11'd997 ) |
 ( (snoop_in == cam_loc998[14:0]) ? cam_loc998 : 11'd998 ) |
 ( (snoop_in == cam_loc999[14:0]) ? cam_loc999 : 11'd999 ) |
 ( (snoop_in == cam_loc1000[14:0]) ? cam_loc1000 : 11'd1000 ) |
 ( (snoop_in == cam_loc1001[14:0]) ? cam_loc1001 : 11'd1001 ) |
 ( (snoop_in == cam_loc1002[14:0]) ? cam_loc1002 : 11'd1002 ) |
 ( (snoop_in == cam_loc1003[14:0]) ? cam_loc1003 : 11'd1003 ) |
 ( (snoop_in == cam_loc1004[14:0]) ? cam_loc1004 : 11'd1004 ) |
 ( (snoop_in == cam_loc1005[14:0]) ? cam_loc1005 : 11'd1005 ) |
 ( (snoop_in == cam_loc1006[14:0]) ? cam_loc1006 : 11'd1006 ) |
 ( (snoop_in == cam_loc1007[14:0]) ? cam_loc1007 : 11'd1007 ) |
 ( (snoop_in == cam_loc1008[14:0]) ? cam_loc1008 : 11'd1008 ) |
 ( (snoop_in == cam_loc1009[14:0]) ? cam_loc1009 : 11'd1009 ) |
 ( (snoop_in == cam_loc1010[14:0]) ? cam_loc1010 : 11'd1010 ) |
 ( (snoop_in == cam_loc1011[14:0]) ? cam_loc1011 : 11'd1011 ) |
 ( (snoop_in == cam_loc1012[14:0]) ? cam_loc1012 : 11'd1012 ) |
 ( (snoop_in == cam_loc1013[14:0]) ? cam_loc1013 : 11'd1013 ) |
 ( (snoop_in == cam_loc1014[14:0]) ? cam_loc1014 : 11'd1014 ) |
 ( (snoop_in == cam_loc1015[14:0]) ? cam_loc1015 : 11'd1015 ) |
 ( (snoop_in == cam_loc1016[14:0]) ? cam_loc1016 : 11'd1016 ) |
 ( (snoop_in == cam_loc1017[14:0]) ? cam_loc1017 : 11'd1017 ) |
 ( (snoop_in == cam_loc1018[14:0]) ? cam_loc1018 : 11'd1018 ) |
 ( (snoop_in == cam_loc1019[14:0]) ? cam_loc1019 : 11'd1019 ) |
 ( (snoop_in == cam_loc1020[14:0]) ? cam_loc1020 : 11'd1020 ) |
 ( (snoop_in == cam_loc1021[14:0]) ? cam_loc1021 : 11'd1021 ) |
 ( (snoop_in == cam_loc1022[14:0]) ? cam_loc1022 : 11'd1022 ) |
 ( (snoop_in == cam_loc1023[14:0]) ? cam_loc1023 : 11'd1023 ) |
 ( (snoop_in == cam_loc1024[14:0]) ? cam_loc1024 : 11'd1024 ) |
 ( (snoop_in == cam_loc1025[14:0]) ? cam_loc1025 : 11'd1025 ) |
 ( (snoop_in == cam_loc1026[14:0]) ? cam_loc1026 : 11'd1026 ) |
 ( (snoop_in == cam_loc1027[14:0]) ? cam_loc1027 : 11'd1027 ) |
 ( (snoop_in == cam_loc1028[14:0]) ? cam_loc1028 : 11'd1028 ) |
 ( (snoop_in == cam_loc1029[14:0]) ? cam_loc1029 : 11'd1029 ) |
 ( (snoop_in == cam_loc1030[14:0]) ? cam_loc1030 : 11'd1030 ) |
 ( (snoop_in == cam_loc1031[14:0]) ? cam_loc1031 : 11'd1031 ) |
 ( (snoop_in == cam_loc1032[14:0]) ? cam_loc1032 : 11'd1032 ) |
 ( (snoop_in == cam_loc1033[14:0]) ? cam_loc1033 : 11'd1033 ) |
 ( (snoop_in == cam_loc1034[14:0]) ? cam_loc1034 : 11'd1034 ) |
 ( (snoop_in == cam_loc1035[14:0]) ? cam_loc1035 : 11'd1035 ) |
 ( (snoop_in == cam_loc1036[14:0]) ? cam_loc1036 : 11'd1036 ) |
 ( (snoop_in == cam_loc1037[14:0]) ? cam_loc1037 : 11'd1037 ) |
 ( (snoop_in == cam_loc1038[14:0]) ? cam_loc1038 : 11'd1038 ) |
 ( (snoop_in == cam_loc1039[14:0]) ? cam_loc1039 : 11'd1039 ) |
 ( (snoop_in == cam_loc1040[14:0]) ? cam_loc1040 : 11'd1040 ) |
 ( (snoop_in == cam_loc1041[14:0]) ? cam_loc1041 : 11'd1041 ) |
 ( (snoop_in == cam_loc1042[14:0]) ? cam_loc1042 : 11'd1042 ) |
 ( (snoop_in == cam_loc1043[14:0]) ? cam_loc1043 : 11'd1043 ) |
 ( (snoop_in == cam_loc1044[14:0]) ? cam_loc1044 : 11'd1044 ) |
 ( (snoop_in == cam_loc1045[14:0]) ? cam_loc1045 : 11'd1045 ) |
 ( (snoop_in == cam_loc1046[14:0]) ? cam_loc1046 : 11'd1046 ) |
 ( (snoop_in == cam_loc1047[14:0]) ? cam_loc1047 : 11'd1047 ) |
 ( (snoop_in == cam_loc1048[14:0]) ? cam_loc1048 : 11'd1048 ) |
 ( (snoop_in == cam_loc1049[14:0]) ? cam_loc1049 : 11'd1049 ) |
 ( (snoop_in == cam_loc1050[14:0]) ? cam_loc1050 : 11'd1050 ) |
 ( (snoop_in == cam_loc1051[14:0]) ? cam_loc1051 : 11'd1051 ) |
 ( (snoop_in == cam_loc1052[14:0]) ? cam_loc1052 : 11'd1052 ) |
 ( (snoop_in == cam_loc1053[14:0]) ? cam_loc1053 : 11'd1053 ) |
 ( (snoop_in == cam_loc1054[14:0]) ? cam_loc1054 : 11'd1054 ) |
 ( (snoop_in == cam_loc1055[14:0]) ? cam_loc1055 : 11'd1055 ) |
 ( (snoop_in == cam_loc1056[14:0]) ? cam_loc1056 : 11'd1056 ) |
 ( (snoop_in == cam_loc1057[14:0]) ? cam_loc1057 : 11'd1057 ) |
 ( (snoop_in == cam_loc1058[14:0]) ? cam_loc1058 : 11'd1058 ) |
 ( (snoop_in == cam_loc1059[14:0]) ? cam_loc1059 : 11'd1059 ) |
 ( (snoop_in == cam_loc1060[14:0]) ? cam_loc1060 : 11'd1060 ) |
 ( (snoop_in == cam_loc1061[14:0]) ? cam_loc1061 : 11'd1061 ) |
 ( (snoop_in == cam_loc1062[14:0]) ? cam_loc1062 : 11'd1062 ) |
 ( (snoop_in == cam_loc1063[14:0]) ? cam_loc1063 : 11'd1063 ) |
 ( (snoop_in == cam_loc1064[14:0]) ? cam_loc1064 : 11'd1064 ) |
 ( (snoop_in == cam_loc1065[14:0]) ? cam_loc1065 : 11'd1065 ) |
 ( (snoop_in == cam_loc1066[14:0]) ? cam_loc1066 : 11'd1066 ) |
 ( (snoop_in == cam_loc1067[14:0]) ? cam_loc1067 : 11'd1067 ) |
 ( (snoop_in == cam_loc1068[14:0]) ? cam_loc1068 : 11'd1068 ) |
 ( (snoop_in == cam_loc1069[14:0]) ? cam_loc1069 : 11'd1069 ) |
 ( (snoop_in == cam_loc1070[14:0]) ? cam_loc1070 : 11'd1070 ) |
 ( (snoop_in == cam_loc1071[14:0]) ? cam_loc1071 : 11'd1071 ) |
 ( (snoop_in == cam_loc1072[14:0]) ? cam_loc1072 : 11'd1072 ) |
 ( (snoop_in == cam_loc1073[14:0]) ? cam_loc1073 : 11'd1073 ) |
 ( (snoop_in == cam_loc1074[14:0]) ? cam_loc1074 : 11'd1074 ) |
 ( (snoop_in == cam_loc1075[14:0]) ? cam_loc1075 : 11'd1075 ) |
 ( (snoop_in == cam_loc1076[14:0]) ? cam_loc1076 : 11'd1076 ) |
 ( (snoop_in == cam_loc1077[14:0]) ? cam_loc1077 : 11'd1077 ) |
 ( (snoop_in == cam_loc1078[14:0]) ? cam_loc1078 : 11'd1078 ) |
 ( (snoop_in == cam_loc1079[14:0]) ? cam_loc1079 : 11'd1079 ) |
 ( (snoop_in == cam_loc1080[14:0]) ? cam_loc1080 : 11'd1080 ) |
 ( (snoop_in == cam_loc1081[14:0]) ? cam_loc1081 : 11'd1081 ) |
 ( (snoop_in == cam_loc1082[14:0]) ? cam_loc1082 : 11'd1082 ) |
 ( (snoop_in == cam_loc1083[14:0]) ? cam_loc1083 : 11'd1083 ) |
 ( (snoop_in == cam_loc1084[14:0]) ? cam_loc1084 : 11'd1084 ) |
 ( (snoop_in == cam_loc1085[14:0]) ? cam_loc1085 : 11'd1085 ) |
 ( (snoop_in == cam_loc1086[14:0]) ? cam_loc1086 : 11'd1086 ) |
 ( (snoop_in == cam_loc1087[14:0]) ? cam_loc1087 : 11'd1087 ) |
 ( (snoop_in == cam_loc1088[14:0]) ? cam_loc1088 : 11'd1088 ) |
 ( (snoop_in == cam_loc1089[14:0]) ? cam_loc1089 : 11'd1089 ) |
 ( (snoop_in == cam_loc1090[14:0]) ? cam_loc1090 : 11'd1090 ) |
 ( (snoop_in == cam_loc1091[14:0]) ? cam_loc1091 : 11'd1091 ) |
 ( (snoop_in == cam_loc1092[14:0]) ? cam_loc1092 : 11'd1092 ) |
 ( (snoop_in == cam_loc1093[14:0]) ? cam_loc1093 : 11'd1093 ) |
 ( (snoop_in == cam_loc1094[14:0]) ? cam_loc1094 : 11'd1094 ) |
 ( (snoop_in == cam_loc1095[14:0]) ? cam_loc1095 : 11'd1095 ) |
 ( (snoop_in == cam_loc1096[14:0]) ? cam_loc1096 : 11'd1096 ) |
 ( (snoop_in == cam_loc1097[14:0]) ? cam_loc1097 : 11'd1097 ) |
 ( (snoop_in == cam_loc1098[14:0]) ? cam_loc1098 : 11'd1098 ) |
 ( (snoop_in == cam_loc1099[14:0]) ? cam_loc1099 : 11'd1099 )

;

wire assign freedup_loc_valid = snoop_match;

endmodule
